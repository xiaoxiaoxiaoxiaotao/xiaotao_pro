`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2020/08/18 21:58:31
// Design Name: 
// Module Name: sparse_mxv_top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

`define counter 1024
`define newcounter 1031
module sparse_mxv_top(
    input clk,
    input rst,
    input idle,
    input [1023:0] inputx_output,
    input [1023:0] inputw0,
   input [1023:0] inputw1,

   input [1023:0] inputw4,
   input [1023:0] inputw5,

   input [1023:0] inputw8,
   input [1023:0] inputw9,

   input [1023:0] inputw12,
   input [1023:0] inputw13,

    input [159:0] inputw0_index,
   input [159:0] inputw1_index,

   input [159:0] inputw4_index,
   input [159:0] inputw5_index,

   input [159:0] inputw8_index,
   input [159:0] inputw9_index,

   input [159:0] inputw12_index,
   input [159:0] inputw13_index,


    output reg [15:0] one_elements,
    output reg [15:0] one_elements1,

    output reg [15:0] one_elements4,
    output reg [15:0] one_elements5,

    output reg [15:0] one_elements8,
    output reg [15:0] one_elements9,

    output reg [15:0] one_elements12,
    output reg [15:0] one_elements13

    );
// the module of sparse matrix X  dence vector 
// latency is 30
    // reg to store temp result
    reg  [511:0]   active_xt       [31:0] ;


  
    wire [15:0]    temp0_result_32  [31:0];
    reg  [15:0]    temp0_result_16  [15:0];
    reg  [15:0]    temp0_result_8   [7:0];
    reg  [15:0]    temp0_result_4   [3:0];
    reg  [15:0]    temp0_result_2   [1:0]; 


    wire [15:0]    temp1_result_32  [31:0];
    reg  [15:0]    temp1_result_16  [15:0];
    reg  [15:0]    temp1_result_8   [7:0];
    reg  [15:0]    temp1_result_4   [3:0];
    reg  [15:0]    temp1_result_2   [1:0]; 


   

    wire [15:0]    temp4_result_32  [31:0];
    reg  [15:0]    temp4_result_16  [15:0];
    reg  [15:0]    temp4_result_8   [7:0];
    reg  [15:0]    temp4_result_4   [3:0];
    reg  [15:0]    temp4_result_2   [1:0]; 


    wire [15:0]    temp5_result_32  [31:0];
    reg  [15:0]    temp5_result_16  [15:0];
    reg  [15:0]    temp5_result_8   [7:0];
    reg  [15:0]    temp5_result_4   [3:0];
    reg  [15:0]    temp5_result_2   [1:0]; 


   

    wire [15:0]    temp8_result_32  [31:0];
    reg  [15:0]    temp8_result_16  [15:0];
    reg  [15:0]    temp8_result_8   [7:0];
    reg  [15:0]    temp8_result_4   [3:0];
    reg  [15:0]    temp8_result_2   [1:0]; 


    wire [15:0]    temp9_result_32  [31:0];
    reg  [15:0]    temp9_result_16  [15:0];
    reg  [15:0]    temp9_result_8   [7:0];
    reg  [15:0]    temp9_result_4   [3:0];
    reg  [15:0]    temp9_result_2   [1:0]; 


   

    wire [15:0]    temp12_result_32  [31:0];
    reg  [15:0]    temp12_result_16  [15:0];
    reg  [15:0]    temp12_result_8   [7:0];
    reg  [15:0]    temp12_result_4   [3:0];
    reg  [15:0]    temp12_result_2   [1:0]; 


    wire [15:0]    temp13_result_32  [31:0];
    reg  [15:0]    temp13_result_16  [15:0];
    reg  [15:0]    temp13_result_8   [7:0];
    reg  [15:0]    temp13_result_4   [3:0];
    reg  [15:0]    temp13_result_2   [1:0]; 


    //control signal 
    
    reg    spmvidle ;
    reg    spmvidle1;
    reg    spmvidle2;
    reg    spmvidle3;

    
    reg    [4:0] state ;
    reg    [31:0] statecount ;


    // state parameter
    parameter  Start                                                       =    0;
    parameter  Load0                                                       =    27;
    parameter  Load1                                                       =    1;
    parameter  Load2                                                       =    2;
    parameter  Load3                                                       =    3;
    parameter  Load4                                                       =    25;
    parameter  Wait1                                                       =    4;
    parameter  Wait2                                                       =    5;
    parameter  Wait3                                                       =    6;
    parameter  Wait4                                                       =    7;
    parameter  Wait5                                                       =    8;
    parameter  Wait6                                                       =    9;
    parameter  Wait7                                                       =    26;
    parameter  Wait_Add128to64                                             =    10;
    parameter  Wait_Add128to64_64to32                                      =    11;
    parameter  Wait_Add128to64_64to32_32to16                               =    12;
    parameter  Wait_Add128to64_64to32_32to16_16to8                         =    13;
    parameter  Wait_Add128to64_64to32_32to16_16to8_8to4                    =    14;
    parameter  Wait_Add128to64_64to32_32to16_16to8_8to4_4to2               =    15;
    parameter  Wait_Add128to64_64to32_32to16_16to8_8to4_4to2_2to1          =    16;
    parameter  Add128to64_64to32_32to16_16to8_8to4_4to2_2to1               =    17;
    parameter  Add64to32_32to16_16to8_8to4_4to2_2to1                       =    18;
    parameter  Add32to16_16to8_8to4_4to2_2to1                              =    19;
    parameter  Add16to8_8to4_4to2_2to1                                     =    20;
    parameter  Add8to4_4to2_2to1                                           =    21;
    parameter  Add4to2_2to1                                                =    22;
    parameter  Add2to1                                                     =    23;
    parameter  Stop                                                        =    24;


    

   
sparse_mxv sparse0_mxv0(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[0]),.inputw(inputw0[31:0]),.inputw_index(inputw0_index[19:0]),.counter(`counter),.output_onebank(temp0_result_32[0]));
sparse_mxv sparse0_mxv1(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[1]),.inputw(inputw0[63:32]),.inputw_index(inputw0_index[19:0]),.counter(`counter),.output_onebank(temp0_result_32[1]));
sparse_mxv sparse0_mxv2(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[2]),.inputw(inputw0[95:64]),.inputw_index(inputw0_index[19:0]),.counter(`counter),.output_onebank(temp0_result_32[2]));
sparse_mxv sparse0_mxv3(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[3]),.inputw(inputw0[127:96]),.inputw_index(inputw0_index[19:0]),.counter(`counter),.output_onebank(temp0_result_32[3]));
sparse_mxv sparse0_mxv4(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[4]),.inputw(inputw0[159:128]),.inputw_index(inputw0_index[39:20]),.counter(`counter),.output_onebank(temp0_result_32[4]));
sparse_mxv sparse0_mxv5(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[5]),.inputw(inputw0[191:160]),.inputw_index(inputw0_index[39:20]),.counter(`counter),.output_onebank(temp0_result_32[5]));
sparse_mxv sparse0_mxv6(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[6]),.inputw(inputw0[223:192]),.inputw_index(inputw0_index[39:20]),.counter(`counter),.output_onebank(temp0_result_32[6]));
sparse_mxv sparse0_mxv7(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[7]),.inputw(inputw0[255:224]),.inputw_index(inputw0_index[39:20]),.counter(`counter),.output_onebank(temp0_result_32[7]));
sparse_mxv sparse0_mxv8(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[8]),.inputw(inputw0[287:256]),.inputw_index(inputw0_index[59:40]),.counter(`counter),.output_onebank(temp0_result_32[8]));
sparse_mxv sparse0_mxv9(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[9]),.inputw(inputw0[319:288]),.inputw_index(inputw0_index[59:40]),.counter(`counter),.output_onebank(temp0_result_32[9]));
sparse_mxv sparse0_mxv10(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[10]),.inputw(inputw0[351:320]),.inputw_index(inputw0_index[59:40]),.counter(`counter),.output_onebank(temp0_result_32[10]));
sparse_mxv sparse0_mxv11(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[11]),.inputw(inputw0[383:352]),.inputw_index(inputw0_index[59:40]),.counter(`counter),.output_onebank(temp0_result_32[11]));
sparse_mxv sparse0_mxv12(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[12]),.inputw(inputw0[415:384]),.inputw_index(inputw0_index[79:60]),.counter(`counter),.output_onebank(temp0_result_32[12]));
sparse_mxv sparse0_mxv13(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[13]),.inputw(inputw0[447:416]),.inputw_index(inputw0_index[79:60]),.counter(`counter),.output_onebank(temp0_result_32[13]));
sparse_mxv sparse0_mxv14(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[14]),.inputw(inputw0[479:448]),.inputw_index(inputw0_index[79:60]),.counter(`counter),.output_onebank(temp0_result_32[14]));
sparse_mxv sparse0_mxv15(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[15]),.inputw(inputw0[511:480]),.inputw_index(inputw0_index[79:60]),.counter(`counter),.output_onebank(temp0_result_32[15]));
sparse_mxv sparse0_mxv16(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[16]),.inputw(inputw0[543:512]),.inputw_index(inputw0_index[99:80]),.counter(`counter),.output_onebank(temp0_result_32[16]));
sparse_mxv sparse0_mxv17(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[17]),.inputw(inputw0[575:544]),.inputw_index(inputw0_index[99:80]),.counter(`counter),.output_onebank(temp0_result_32[17]));
sparse_mxv sparse0_mxv18(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[18]),.inputw(inputw0[607:576]),.inputw_index(inputw0_index[99:80]),.counter(`counter),.output_onebank(temp0_result_32[18]));
sparse_mxv sparse0_mxv19(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[19]),.inputw(inputw0[639:608]),.inputw_index(inputw0_index[99:80]),.counter(`counter),.output_onebank(temp0_result_32[19]));
sparse_mxv sparse0_mxv20(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[20]),.inputw(inputw0[671:640]),.inputw_index(inputw0_index[119:100]),.counter(`counter),.output_onebank(temp0_result_32[20]));
sparse_mxv sparse0_mxv21(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[21]),.inputw(inputw0[703:672]),.inputw_index(inputw0_index[119:100]),.counter(`counter),.output_onebank(temp0_result_32[21]));
sparse_mxv sparse0_mxv22(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[22]),.inputw(inputw0[735:704]),.inputw_index(inputw0_index[119:100]),.counter(`counter),.output_onebank(temp0_result_32[22]));
sparse_mxv sparse0_mxv23(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[23]),.inputw(inputw0[767:736]),.inputw_index(inputw0_index[119:100]),.counter(`counter),.output_onebank(temp0_result_32[23]));
sparse_mxv sparse0_mxv24(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[24]),.inputw(inputw0[799:768]),.inputw_index(inputw0_index[139:120]),.counter(`counter),.output_onebank(temp0_result_32[24]));
sparse_mxv sparse0_mxv25(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[25]),.inputw(inputw0[831:800]),.inputw_index(inputw0_index[139:120]),.counter(`counter),.output_onebank(temp0_result_32[25]));
sparse_mxv sparse0_mxv26(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[26]),.inputw(inputw0[863:832]),.inputw_index(inputw0_index[139:120]),.counter(`counter),.output_onebank(temp0_result_32[26]));
sparse_mxv sparse0_mxv27(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[27]),.inputw(inputw0[895:864]),.inputw_index(inputw0_index[139:120]),.counter(`counter),.output_onebank(temp0_result_32[27]));
sparse_mxv sparse0_mxv28(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[28]),.inputw(inputw0[927:896]),.inputw_index(inputw0_index[159:140]),.counter(`counter),.output_onebank(temp0_result_32[28]));
sparse_mxv sparse0_mxv29(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[29]),.inputw(inputw0[959:928]),.inputw_index(inputw0_index[159:140]),.counter(`counter),.output_onebank(temp0_result_32[29]));
sparse_mxv sparse0_mxv30(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[30]),.inputw(inputw0[991:960]),.inputw_index(inputw0_index[159:140]),.counter(`counter),.output_onebank(temp0_result_32[30]));
sparse_mxv sparse0_mxv31(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[31]),.inputw(inputw0[1023:992]),.inputw_index(inputw0_index[159:140]),.counter(`counter),.output_onebank(temp0_result_32[31]));
sparse_mxv sparse1_mxv0(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[0]),.inputw(inputw1[31:0]),.inputw_index(inputw1_index[19:0]),.counter(`counter),.output_onebank(temp1_result_32[0]));
sparse_mxv sparse1_mxv1(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[1]),.inputw(inputw1[63:32]),.inputw_index(inputw1_index[19:0]),.counter(`counter),.output_onebank(temp1_result_32[1]));
sparse_mxv sparse1_mxv2(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[2]),.inputw(inputw1[95:64]),.inputw_index(inputw1_index[19:0]),.counter(`counter),.output_onebank(temp1_result_32[2]));
sparse_mxv sparse1_mxv3(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[3]),.inputw(inputw1[127:96]),.inputw_index(inputw1_index[19:0]),.counter(`counter),.output_onebank(temp1_result_32[3]));
sparse_mxv sparse1_mxv4(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[4]),.inputw(inputw1[159:128]),.inputw_index(inputw1_index[39:20]),.counter(`counter),.output_onebank(temp1_result_32[4]));
sparse_mxv sparse1_mxv5(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[5]),.inputw(inputw1[191:160]),.inputw_index(inputw1_index[39:20]),.counter(`counter),.output_onebank(temp1_result_32[5]));
sparse_mxv sparse1_mxv6(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[6]),.inputw(inputw1[223:192]),.inputw_index(inputw1_index[39:20]),.counter(`counter),.output_onebank(temp1_result_32[6]));
sparse_mxv sparse1_mxv7(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[7]),.inputw(inputw1[255:224]),.inputw_index(inputw1_index[39:20]),.counter(`counter),.output_onebank(temp1_result_32[7]));
sparse_mxv sparse1_mxv8(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[8]),.inputw(inputw1[287:256]),.inputw_index(inputw1_index[59:40]),.counter(`counter),.output_onebank(temp1_result_32[8]));
sparse_mxv sparse1_mxv9(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[9]),.inputw(inputw1[319:288]),.inputw_index(inputw1_index[59:40]),.counter(`counter),.output_onebank(temp1_result_32[9]));
sparse_mxv sparse1_mxv10(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[10]),.inputw(inputw1[351:320]),.inputw_index(inputw1_index[59:40]),.counter(`counter),.output_onebank(temp1_result_32[10]));
sparse_mxv sparse1_mxv11(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[11]),.inputw(inputw1[383:352]),.inputw_index(inputw1_index[59:40]),.counter(`counter),.output_onebank(temp1_result_32[11]));
sparse_mxv sparse1_mxv12(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[12]),.inputw(inputw1[415:384]),.inputw_index(inputw1_index[79:60]),.counter(`counter),.output_onebank(temp1_result_32[12]));
sparse_mxv sparse1_mxv13(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[13]),.inputw(inputw1[447:416]),.inputw_index(inputw1_index[79:60]),.counter(`counter),.output_onebank(temp1_result_32[13]));
sparse_mxv sparse1_mxv14(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[14]),.inputw(inputw1[479:448]),.inputw_index(inputw1_index[79:60]),.counter(`counter),.output_onebank(temp1_result_32[14]));
sparse_mxv sparse1_mxv15(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[15]),.inputw(inputw1[511:480]),.inputw_index(inputw1_index[79:60]),.counter(`counter),.output_onebank(temp1_result_32[15]));
sparse_mxv sparse1_mxv16(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[16]),.inputw(inputw1[543:512]),.inputw_index(inputw1_index[99:80]),.counter(`counter),.output_onebank(temp1_result_32[16]));
sparse_mxv sparse1_mxv17(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[17]),.inputw(inputw1[575:544]),.inputw_index(inputw1_index[99:80]),.counter(`counter),.output_onebank(temp1_result_32[17]));
sparse_mxv sparse1_mxv18(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[18]),.inputw(inputw1[607:576]),.inputw_index(inputw1_index[99:80]),.counter(`counter),.output_onebank(temp1_result_32[18]));
sparse_mxv sparse1_mxv19(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[19]),.inputw(inputw1[639:608]),.inputw_index(inputw1_index[99:80]),.counter(`counter),.output_onebank(temp1_result_32[19]));
sparse_mxv sparse1_mxv20(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[20]),.inputw(inputw1[671:640]),.inputw_index(inputw1_index[119:100]),.counter(`counter),.output_onebank(temp1_result_32[20]));
sparse_mxv sparse1_mxv21(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[21]),.inputw(inputw1[703:672]),.inputw_index(inputw1_index[119:100]),.counter(`counter),.output_onebank(temp1_result_32[21]));
sparse_mxv sparse1_mxv22(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[22]),.inputw(inputw1[735:704]),.inputw_index(inputw1_index[119:100]),.counter(`counter),.output_onebank(temp1_result_32[22]));
sparse_mxv sparse1_mxv23(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[23]),.inputw(inputw1[767:736]),.inputw_index(inputw1_index[119:100]),.counter(`counter),.output_onebank(temp1_result_32[23]));
sparse_mxv sparse1_mxv24(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[24]),.inputw(inputw1[799:768]),.inputw_index(inputw1_index[139:120]),.counter(`counter),.output_onebank(temp1_result_32[24]));
sparse_mxv sparse1_mxv25(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[25]),.inputw(inputw1[831:800]),.inputw_index(inputw1_index[139:120]),.counter(`counter),.output_onebank(temp1_result_32[25]));
sparse_mxv sparse1_mxv26(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[26]),.inputw(inputw1[863:832]),.inputw_index(inputw1_index[139:120]),.counter(`counter),.output_onebank(temp1_result_32[26]));
sparse_mxv sparse1_mxv27(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[27]),.inputw(inputw1[895:864]),.inputw_index(inputw1_index[139:120]),.counter(`counter),.output_onebank(temp1_result_32[27]));
sparse_mxv sparse1_mxv28(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[28]),.inputw(inputw1[927:896]),.inputw_index(inputw1_index[159:140]),.counter(`counter),.output_onebank(temp1_result_32[28]));
sparse_mxv sparse1_mxv29(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[29]),.inputw(inputw1[959:928]),.inputw_index(inputw1_index[159:140]),.counter(`counter),.output_onebank(temp1_result_32[29]));
sparse_mxv sparse1_mxv30(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[30]),.inputw(inputw1[991:960]),.inputw_index(inputw1_index[159:140]),.counter(`counter),.output_onebank(temp1_result_32[30]));
sparse_mxv sparse1_mxv31(.clk(clk),.idle(spmvidle2),.rst(rst),.inputx(active_xt[31]),.inputw(inputw1[1023:992]),.inputw_index(inputw1_index[159:140]),.counter(`counter),.output_onebank(temp1_result_32[31]));


sparse_mxv sparse4_mxv0(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[0]),.inputw(inputw4[31:0]),.inputw_index(inputw4_index[19:0]),.counter(`counter),.output_onebank(temp4_result_32[0]));
sparse_mxv sparse4_mxv1(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[1]),.inputw(inputw4[63:32]),.inputw_index(inputw4_index[19:0]),.counter(`counter),.output_onebank(temp4_result_32[1]));
sparse_mxv sparse4_mxv2(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[2]),.inputw(inputw4[95:64]),.inputw_index(inputw4_index[19:0]),.counter(`counter),.output_onebank(temp4_result_32[2]));
sparse_mxv sparse4_mxv3(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[3]),.inputw(inputw4[127:96]),.inputw_index(inputw4_index[19:0]),.counter(`counter),.output_onebank(temp4_result_32[3]));
sparse_mxv sparse4_mxv4(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[4]),.inputw(inputw4[159:128]),.inputw_index(inputw4_index[39:20]),.counter(`counter),.output_onebank(temp4_result_32[4]));
sparse_mxv sparse4_mxv5(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[5]),.inputw(inputw4[191:160]),.inputw_index(inputw4_index[39:20]),.counter(`counter),.output_onebank(temp4_result_32[5]));
sparse_mxv sparse4_mxv6(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[6]),.inputw(inputw4[223:192]),.inputw_index(inputw4_index[39:20]),.counter(`counter),.output_onebank(temp4_result_32[6]));
sparse_mxv sparse4_mxv7(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[7]),.inputw(inputw4[255:224]),.inputw_index(inputw4_index[39:20]),.counter(`counter),.output_onebank(temp4_result_32[7]));
sparse_mxv sparse4_mxv8(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[8]),.inputw(inputw4[287:256]),.inputw_index(inputw4_index[59:40]),.counter(`counter),.output_onebank(temp4_result_32[8]));
sparse_mxv sparse4_mxv9(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[9]),.inputw(inputw4[319:288]),.inputw_index(inputw4_index[59:40]),.counter(`counter),.output_onebank(temp4_result_32[9]));
sparse_mxv sparse4_mxv10(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[10]),.inputw(inputw4[351:320]),.inputw_index(inputw4_index[59:40]),.counter(`counter),.output_onebank(temp4_result_32[10]));
sparse_mxv sparse4_mxv11(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[11]),.inputw(inputw4[383:352]),.inputw_index(inputw4_index[59:40]),.counter(`counter),.output_onebank(temp4_result_32[11]));
sparse_mxv sparse4_mxv12(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[12]),.inputw(inputw4[415:384]),.inputw_index(inputw4_index[79:60]),.counter(`counter),.output_onebank(temp4_result_32[12]));
sparse_mxv sparse4_mxv13(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[13]),.inputw(inputw4[447:416]),.inputw_index(inputw4_index[79:60]),.counter(`counter),.output_onebank(temp4_result_32[13]));
sparse_mxv sparse4_mxv14(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[14]),.inputw(inputw4[479:448]),.inputw_index(inputw4_index[79:60]),.counter(`counter),.output_onebank(temp4_result_32[14]));
sparse_mxv sparse4_mxv15(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[15]),.inputw(inputw4[511:480]),.inputw_index(inputw4_index[79:60]),.counter(`counter),.output_onebank(temp4_result_32[15]));
sparse_mxv sparse4_mxv16(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[16]),.inputw(inputw4[543:512]),.inputw_index(inputw4_index[99:80]),.counter(`counter),.output_onebank(temp4_result_32[16]));
sparse_mxv sparse4_mxv17(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[17]),.inputw(inputw4[575:544]),.inputw_index(inputw4_index[99:80]),.counter(`counter),.output_onebank(temp4_result_32[17]));
sparse_mxv sparse4_mxv18(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[18]),.inputw(inputw4[607:576]),.inputw_index(inputw4_index[99:80]),.counter(`counter),.output_onebank(temp4_result_32[18]));
sparse_mxv sparse4_mxv19(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[19]),.inputw(inputw4[639:608]),.inputw_index(inputw4_index[99:80]),.counter(`counter),.output_onebank(temp4_result_32[19]));
sparse_mxv sparse4_mxv20(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[20]),.inputw(inputw4[671:640]),.inputw_index(inputw4_index[119:100]),.counter(`counter),.output_onebank(temp4_result_32[20]));
sparse_mxv sparse4_mxv21(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[21]),.inputw(inputw4[703:672]),.inputw_index(inputw4_index[119:100]),.counter(`counter),.output_onebank(temp4_result_32[21]));
sparse_mxv sparse4_mxv22(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[22]),.inputw(inputw4[735:704]),.inputw_index(inputw4_index[119:100]),.counter(`counter),.output_onebank(temp4_result_32[22]));
sparse_mxv sparse4_mxv23(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[23]),.inputw(inputw4[767:736]),.inputw_index(inputw4_index[119:100]),.counter(`counter),.output_onebank(temp4_result_32[23]));
sparse_mxv sparse4_mxv24(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[24]),.inputw(inputw4[799:768]),.inputw_index(inputw4_index[139:120]),.counter(`counter),.output_onebank(temp4_result_32[24]));
sparse_mxv sparse4_mxv25(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[25]),.inputw(inputw4[831:800]),.inputw_index(inputw4_index[139:120]),.counter(`counter),.output_onebank(temp4_result_32[25]));
sparse_mxv sparse4_mxv26(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[26]),.inputw(inputw4[863:832]),.inputw_index(inputw4_index[139:120]),.counter(`counter),.output_onebank(temp4_result_32[26]));
sparse_mxv sparse4_mxv27(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[27]),.inputw(inputw4[895:864]),.inputw_index(inputw4_index[139:120]),.counter(`counter),.output_onebank(temp4_result_32[27]));
sparse_mxv sparse4_mxv28(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[28]),.inputw(inputw4[927:896]),.inputw_index(inputw4_index[159:140]),.counter(`counter),.output_onebank(temp4_result_32[28]));
sparse_mxv sparse4_mxv29(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[29]),.inputw(inputw4[959:928]),.inputw_index(inputw4_index[159:140]),.counter(`counter),.output_onebank(temp4_result_32[29]));
sparse_mxv sparse4_mxv30(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[30]),.inputw(inputw4[991:960]),.inputw_index(inputw4_index[159:140]),.counter(`counter),.output_onebank(temp4_result_32[30]));
sparse_mxv sparse4_mxv31(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[31]),.inputw(inputw4[1023:992]),.inputw_index(inputw4_index[159:140]),.counter(`counter),.output_onebank(temp4_result_32[31]));
sparse_mxv sparse5_mxv0(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[0]),.inputw(inputw5[31:0]),.inputw_index(inputw5_index[19:0]),.counter(`counter),.output_onebank(temp5_result_32[0]));
sparse_mxv sparse5_mxv1(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[1]),.inputw(inputw5[63:32]),.inputw_index(inputw5_index[19:0]),.counter(`counter),.output_onebank(temp5_result_32[1]));
sparse_mxv sparse5_mxv2(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[2]),.inputw(inputw5[95:64]),.inputw_index(inputw5_index[19:0]),.counter(`counter),.output_onebank(temp5_result_32[2]));
sparse_mxv sparse5_mxv3(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[3]),.inputw(inputw5[127:96]),.inputw_index(inputw5_index[19:0]),.counter(`counter),.output_onebank(temp5_result_32[3]));
sparse_mxv sparse5_mxv4(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[4]),.inputw(inputw5[159:128]),.inputw_index(inputw5_index[39:20]),.counter(`counter),.output_onebank(temp5_result_32[4]));
sparse_mxv sparse5_mxv5(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[5]),.inputw(inputw5[191:160]),.inputw_index(inputw5_index[39:20]),.counter(`counter),.output_onebank(temp5_result_32[5]));
sparse_mxv sparse5_mxv6(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[6]),.inputw(inputw5[223:192]),.inputw_index(inputw5_index[39:20]),.counter(`counter),.output_onebank(temp5_result_32[6]));
sparse_mxv sparse5_mxv7(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[7]),.inputw(inputw5[255:224]),.inputw_index(inputw5_index[39:20]),.counter(`counter),.output_onebank(temp5_result_32[7]));
sparse_mxv sparse5_mxv8(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[8]),.inputw(inputw5[287:256]),.inputw_index(inputw5_index[59:40]),.counter(`counter),.output_onebank(temp5_result_32[8]));
sparse_mxv sparse5_mxv9(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[9]),.inputw(inputw5[319:288]),.inputw_index(inputw5_index[59:40]),.counter(`counter),.output_onebank(temp5_result_32[9]));
sparse_mxv sparse5_mxv10(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[10]),.inputw(inputw5[351:320]),.inputw_index(inputw5_index[59:40]),.counter(`counter),.output_onebank(temp5_result_32[10]));
sparse_mxv sparse5_mxv11(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[11]),.inputw(inputw5[383:352]),.inputw_index(inputw5_index[59:40]),.counter(`counter),.output_onebank(temp5_result_32[11]));
sparse_mxv sparse5_mxv12(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[12]),.inputw(inputw5[415:384]),.inputw_index(inputw5_index[79:60]),.counter(`counter),.output_onebank(temp5_result_32[12]));
sparse_mxv sparse5_mxv13(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[13]),.inputw(inputw5[447:416]),.inputw_index(inputw5_index[79:60]),.counter(`counter),.output_onebank(temp5_result_32[13]));
sparse_mxv sparse5_mxv14(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[14]),.inputw(inputw5[479:448]),.inputw_index(inputw5_index[79:60]),.counter(`counter),.output_onebank(temp5_result_32[14]));
sparse_mxv sparse5_mxv15(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[15]),.inputw(inputw5[511:480]),.inputw_index(inputw5_index[79:60]),.counter(`counter),.output_onebank(temp5_result_32[15]));
sparse_mxv sparse5_mxv16(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[16]),.inputw(inputw5[543:512]),.inputw_index(inputw5_index[99:80]),.counter(`counter),.output_onebank(temp5_result_32[16]));
sparse_mxv sparse5_mxv17(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[17]),.inputw(inputw5[575:544]),.inputw_index(inputw5_index[99:80]),.counter(`counter),.output_onebank(temp5_result_32[17]));
sparse_mxv sparse5_mxv18(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[18]),.inputw(inputw5[607:576]),.inputw_index(inputw5_index[99:80]),.counter(`counter),.output_onebank(temp5_result_32[18]));
sparse_mxv sparse5_mxv19(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[19]),.inputw(inputw5[639:608]),.inputw_index(inputw5_index[99:80]),.counter(`counter),.output_onebank(temp5_result_32[19]));
sparse_mxv sparse5_mxv20(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[20]),.inputw(inputw5[671:640]),.inputw_index(inputw5_index[119:100]),.counter(`counter),.output_onebank(temp5_result_32[20]));
sparse_mxv sparse5_mxv21(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[21]),.inputw(inputw5[703:672]),.inputw_index(inputw5_index[119:100]),.counter(`counter),.output_onebank(temp5_result_32[21]));
sparse_mxv sparse5_mxv22(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[22]),.inputw(inputw5[735:704]),.inputw_index(inputw5_index[119:100]),.counter(`counter),.output_onebank(temp5_result_32[22]));
sparse_mxv sparse5_mxv23(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[23]),.inputw(inputw5[767:736]),.inputw_index(inputw5_index[119:100]),.counter(`counter),.output_onebank(temp5_result_32[23]));
sparse_mxv sparse5_mxv24(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[24]),.inputw(inputw5[799:768]),.inputw_index(inputw5_index[139:120]),.counter(`counter),.output_onebank(temp5_result_32[24]));
sparse_mxv sparse5_mxv25(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[25]),.inputw(inputw5[831:800]),.inputw_index(inputw5_index[139:120]),.counter(`counter),.output_onebank(temp5_result_32[25]));
sparse_mxv sparse5_mxv26(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[26]),.inputw(inputw5[863:832]),.inputw_index(inputw5_index[139:120]),.counter(`counter),.output_onebank(temp5_result_32[26]));
sparse_mxv sparse5_mxv27(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[27]),.inputw(inputw5[895:864]),.inputw_index(inputw5_index[139:120]),.counter(`counter),.output_onebank(temp5_result_32[27]));
sparse_mxv sparse5_mxv28(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[28]),.inputw(inputw5[927:896]),.inputw_index(inputw5_index[159:140]),.counter(`counter),.output_onebank(temp5_result_32[28]));
sparse_mxv sparse5_mxv29(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[29]),.inputw(inputw5[959:928]),.inputw_index(inputw5_index[159:140]),.counter(`counter),.output_onebank(temp5_result_32[29]));
sparse_mxv sparse5_mxv30(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[30]),.inputw(inputw5[991:960]),.inputw_index(inputw5_index[159:140]),.counter(`counter),.output_onebank(temp5_result_32[30]));
sparse_mxv sparse5_mxv31(.clk(clk),.idle(spmvidle),.rst(rst),.inputx(active_xt[31]),.inputw(inputw5[1023:992]),.inputw_index(inputw5_index[159:140]),.counter(`counter),.output_onebank(temp5_result_32[31]));


sparse_mxv sparse8_mxv0(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[0]),.inputw(inputw8[31:0]),.inputw_index(inputw8_index[19:0]),.counter(`counter),.output_onebank(temp8_result_32[0]));
sparse_mxv sparse8_mxv1(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[1]),.inputw(inputw8[63:32]),.inputw_index(inputw8_index[19:0]),.counter(`counter),.output_onebank(temp8_result_32[1]));
sparse_mxv sparse8_mxv2(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[2]),.inputw(inputw8[95:64]),.inputw_index(inputw8_index[19:0]),.counter(`counter),.output_onebank(temp8_result_32[2]));
sparse_mxv sparse8_mxv3(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[3]),.inputw(inputw8[127:96]),.inputw_index(inputw8_index[19:0]),.counter(`counter),.output_onebank(temp8_result_32[3]));
sparse_mxv sparse8_mxv4(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[4]),.inputw(inputw8[159:128]),.inputw_index(inputw8_index[39:20]),.counter(`counter),.output_onebank(temp8_result_32[4]));
sparse_mxv sparse8_mxv5(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[5]),.inputw(inputw8[191:160]),.inputw_index(inputw8_index[39:20]),.counter(`counter),.output_onebank(temp8_result_32[5]));
sparse_mxv sparse8_mxv6(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[6]),.inputw(inputw8[223:192]),.inputw_index(inputw8_index[39:20]),.counter(`counter),.output_onebank(temp8_result_32[6]));
sparse_mxv sparse8_mxv7(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[7]),.inputw(inputw8[255:224]),.inputw_index(inputw8_index[39:20]),.counter(`counter),.output_onebank(temp8_result_32[7]));
sparse_mxv sparse8_mxv8(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[8]),.inputw(inputw8[287:256]),.inputw_index(inputw8_index[59:40]),.counter(`counter),.output_onebank(temp8_result_32[8]));
sparse_mxv sparse8_mxv9(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[9]),.inputw(inputw8[319:288]),.inputw_index(inputw8_index[59:40]),.counter(`counter),.output_onebank(temp8_result_32[9]));
sparse_mxv sparse8_mxv10(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[10]),.inputw(inputw8[351:320]),.inputw_index(inputw8_index[59:40]),.counter(`counter),.output_onebank(temp8_result_32[10]));
sparse_mxv sparse8_mxv11(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[11]),.inputw(inputw8[383:352]),.inputw_index(inputw8_index[59:40]),.counter(`counter),.output_onebank(temp8_result_32[11]));
sparse_mxv sparse8_mxv12(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[12]),.inputw(inputw8[415:384]),.inputw_index(inputw8_index[79:60]),.counter(`counter),.output_onebank(temp8_result_32[12]));
sparse_mxv sparse8_mxv13(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[13]),.inputw(inputw8[447:416]),.inputw_index(inputw8_index[79:60]),.counter(`counter),.output_onebank(temp8_result_32[13]));
sparse_mxv sparse8_mxv14(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[14]),.inputw(inputw8[479:448]),.inputw_index(inputw8_index[79:60]),.counter(`counter),.output_onebank(temp8_result_32[14]));
sparse_mxv sparse8_mxv15(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[15]),.inputw(inputw8[511:480]),.inputw_index(inputw8_index[79:60]),.counter(`counter),.output_onebank(temp8_result_32[15]));
sparse_mxv sparse8_mxv16(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[16]),.inputw(inputw8[543:512]),.inputw_index(inputw8_index[99:80]),.counter(`counter),.output_onebank(temp8_result_32[16]));
sparse_mxv sparse8_mxv17(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[17]),.inputw(inputw8[575:544]),.inputw_index(inputw8_index[99:80]),.counter(`counter),.output_onebank(temp8_result_32[17]));
sparse_mxv sparse8_mxv18(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[18]),.inputw(inputw8[607:576]),.inputw_index(inputw8_index[99:80]),.counter(`counter),.output_onebank(temp8_result_32[18]));
sparse_mxv sparse8_mxv19(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[19]),.inputw(inputw8[639:608]),.inputw_index(inputw8_index[99:80]),.counter(`counter),.output_onebank(temp8_result_32[19]));
sparse_mxv sparse8_mxv20(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[20]),.inputw(inputw8[671:640]),.inputw_index(inputw8_index[119:100]),.counter(`counter),.output_onebank(temp8_result_32[20]));
sparse_mxv sparse8_mxv21(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[21]),.inputw(inputw8[703:672]),.inputw_index(inputw8_index[119:100]),.counter(`counter),.output_onebank(temp8_result_32[21]));
sparse_mxv sparse8_mxv22(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[22]),.inputw(inputw8[735:704]),.inputw_index(inputw8_index[119:100]),.counter(`counter),.output_onebank(temp8_result_32[22]));
sparse_mxv sparse8_mxv23(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[23]),.inputw(inputw8[767:736]),.inputw_index(inputw8_index[119:100]),.counter(`counter),.output_onebank(temp8_result_32[23]));
sparse_mxv sparse8_mxv24(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[24]),.inputw(inputw8[799:768]),.inputw_index(inputw8_index[139:120]),.counter(`counter),.output_onebank(temp8_result_32[24]));
sparse_mxv sparse8_mxv25(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[25]),.inputw(inputw8[831:800]),.inputw_index(inputw8_index[139:120]),.counter(`counter),.output_onebank(temp8_result_32[25]));
sparse_mxv sparse8_mxv26(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[26]),.inputw(inputw8[863:832]),.inputw_index(inputw8_index[139:120]),.counter(`counter),.output_onebank(temp8_result_32[26]));
sparse_mxv sparse8_mxv27(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[27]),.inputw(inputw8[895:864]),.inputw_index(inputw8_index[139:120]),.counter(`counter),.output_onebank(temp8_result_32[27]));
sparse_mxv sparse8_mxv28(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[28]),.inputw(inputw8[927:896]),.inputw_index(inputw8_index[159:140]),.counter(`counter),.output_onebank(temp8_result_32[28]));
sparse_mxv sparse8_mxv29(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[29]),.inputw(inputw8[959:928]),.inputw_index(inputw8_index[159:140]),.counter(`counter),.output_onebank(temp8_result_32[29]));
sparse_mxv sparse8_mxv30(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[30]),.inputw(inputw8[991:960]),.inputw_index(inputw8_index[159:140]),.counter(`counter),.output_onebank(temp8_result_32[30]));
sparse_mxv sparse8_mxv31(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[31]),.inputw(inputw8[1023:992]),.inputw_index(inputw8_index[159:140]),.counter(`counter),.output_onebank(temp8_result_32[31]));
sparse_mxv sparse9_mxv0(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[0]),.inputw(inputw9[31:0]),.inputw_index(inputw9_index[19:0]),.counter(`counter),.output_onebank(temp9_result_32[0]));
sparse_mxv sparse9_mxv1(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[1]),.inputw(inputw9[63:32]),.inputw_index(inputw9_index[19:0]),.counter(`counter),.output_onebank(temp9_result_32[1]));
sparse_mxv sparse9_mxv2(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[2]),.inputw(inputw9[95:64]),.inputw_index(inputw9_index[19:0]),.counter(`counter),.output_onebank(temp9_result_32[2]));
sparse_mxv sparse9_mxv3(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[3]),.inputw(inputw9[127:96]),.inputw_index(inputw9_index[19:0]),.counter(`counter),.output_onebank(temp9_result_32[3]));
sparse_mxv sparse9_mxv4(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[4]),.inputw(inputw9[159:128]),.inputw_index(inputw9_index[39:20]),.counter(`counter),.output_onebank(temp9_result_32[4]));
sparse_mxv sparse9_mxv5(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[5]),.inputw(inputw9[191:160]),.inputw_index(inputw9_index[39:20]),.counter(`counter),.output_onebank(temp9_result_32[5]));
sparse_mxv sparse9_mxv6(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[6]),.inputw(inputw9[223:192]),.inputw_index(inputw9_index[39:20]),.counter(`counter),.output_onebank(temp9_result_32[6]));
sparse_mxv sparse9_mxv7(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[7]),.inputw(inputw9[255:224]),.inputw_index(inputw9_index[39:20]),.counter(`counter),.output_onebank(temp9_result_32[7]));
sparse_mxv sparse9_mxv8(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[8]),.inputw(inputw9[287:256]),.inputw_index(inputw9_index[59:40]),.counter(`counter),.output_onebank(temp9_result_32[8]));
sparse_mxv sparse9_mxv9(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[9]),.inputw(inputw9[319:288]),.inputw_index(inputw9_index[59:40]),.counter(`counter),.output_onebank(temp9_result_32[9]));
sparse_mxv sparse9_mxv10(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[10]),.inputw(inputw9[351:320]),.inputw_index(inputw9_index[59:40]),.counter(`counter),.output_onebank(temp9_result_32[10]));
sparse_mxv sparse9_mxv11(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[11]),.inputw(inputw9[383:352]),.inputw_index(inputw9_index[59:40]),.counter(`counter),.output_onebank(temp9_result_32[11]));
sparse_mxv sparse9_mxv12(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[12]),.inputw(inputw9[415:384]),.inputw_index(inputw9_index[79:60]),.counter(`counter),.output_onebank(temp9_result_32[12]));
sparse_mxv sparse9_mxv13(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[13]),.inputw(inputw9[447:416]),.inputw_index(inputw9_index[79:60]),.counter(`counter),.output_onebank(temp9_result_32[13]));
sparse_mxv sparse9_mxv14(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[14]),.inputw(inputw9[479:448]),.inputw_index(inputw9_index[79:60]),.counter(`counter),.output_onebank(temp9_result_32[14]));
sparse_mxv sparse9_mxv15(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[15]),.inputw(inputw9[511:480]),.inputw_index(inputw9_index[79:60]),.counter(`counter),.output_onebank(temp9_result_32[15]));
sparse_mxv sparse9_mxv16(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[16]),.inputw(inputw9[543:512]),.inputw_index(inputw9_index[99:80]),.counter(`counter),.output_onebank(temp9_result_32[16]));
sparse_mxv sparse9_mxv17(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[17]),.inputw(inputw9[575:544]),.inputw_index(inputw9_index[99:80]),.counter(`counter),.output_onebank(temp9_result_32[17]));
sparse_mxv sparse9_mxv18(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[18]),.inputw(inputw9[607:576]),.inputw_index(inputw9_index[99:80]),.counter(`counter),.output_onebank(temp9_result_32[18]));
sparse_mxv sparse9_mxv19(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[19]),.inputw(inputw9[639:608]),.inputw_index(inputw9_index[99:80]),.counter(`counter),.output_onebank(temp9_result_32[19]));
sparse_mxv sparse9_mxv20(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[20]),.inputw(inputw9[671:640]),.inputw_index(inputw9_index[119:100]),.counter(`counter),.output_onebank(temp9_result_32[20]));
sparse_mxv sparse9_mxv21(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[21]),.inputw(inputw9[703:672]),.inputw_index(inputw9_index[119:100]),.counter(`counter),.output_onebank(temp9_result_32[21]));
sparse_mxv sparse9_mxv22(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[22]),.inputw(inputw9[735:704]),.inputw_index(inputw9_index[119:100]),.counter(`counter),.output_onebank(temp9_result_32[22]));
sparse_mxv sparse9_mxv23(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[23]),.inputw(inputw9[767:736]),.inputw_index(inputw9_index[119:100]),.counter(`counter),.output_onebank(temp9_result_32[23]));
sparse_mxv sparse9_mxv24(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[24]),.inputw(inputw9[799:768]),.inputw_index(inputw9_index[139:120]),.counter(`counter),.output_onebank(temp9_result_32[24]));
sparse_mxv sparse9_mxv25(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[25]),.inputw(inputw9[831:800]),.inputw_index(inputw9_index[139:120]),.counter(`counter),.output_onebank(temp9_result_32[25]));
sparse_mxv sparse9_mxv26(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[26]),.inputw(inputw9[863:832]),.inputw_index(inputw9_index[139:120]),.counter(`counter),.output_onebank(temp9_result_32[26]));
sparse_mxv sparse9_mxv27(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[27]),.inputw(inputw9[895:864]),.inputw_index(inputw9_index[139:120]),.counter(`counter),.output_onebank(temp9_result_32[27]));
sparse_mxv sparse9_mxv28(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[28]),.inputw(inputw9[927:896]),.inputw_index(inputw9_index[159:140]),.counter(`counter),.output_onebank(temp9_result_32[28]));
sparse_mxv sparse9_mxv29(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[29]),.inputw(inputw9[959:928]),.inputw_index(inputw9_index[159:140]),.counter(`counter),.output_onebank(temp9_result_32[29]));
sparse_mxv sparse9_mxv30(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[30]),.inputw(inputw9[991:960]),.inputw_index(inputw9_index[159:140]),.counter(`counter),.output_onebank(temp9_result_32[30]));
sparse_mxv sparse9_mxv31(.clk(clk),.idle(spmvidle1),.rst(rst),.inputx(active_xt[31]),.inputw(inputw9[1023:992]),.inputw_index(inputw9_index[159:140]),.counter(`counter),.output_onebank(temp9_result_32[31]));


sparse_mxv sparse12_mxv0(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[0]),.inputw(inputw12[31:0]),.inputw_index(inputw12_index[19:0]),.counter(`counter),.output_onebank(temp12_result_32[0]));
sparse_mxv sparse12_mxv1(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[1]),.inputw(inputw12[63:32]),.inputw_index(inputw12_index[19:0]),.counter(`counter),.output_onebank(temp12_result_32[1]));
sparse_mxv sparse12_mxv2(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[2]),.inputw(inputw12[95:64]),.inputw_index(inputw12_index[19:0]),.counter(`counter),.output_onebank(temp12_result_32[2]));
sparse_mxv sparse12_mxv3(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[3]),.inputw(inputw12[127:96]),.inputw_index(inputw12_index[19:0]),.counter(`counter),.output_onebank(temp12_result_32[3]));
sparse_mxv sparse12_mxv4(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[4]),.inputw(inputw12[159:128]),.inputw_index(inputw12_index[39:20]),.counter(`counter),.output_onebank(temp12_result_32[4]));
sparse_mxv sparse12_mxv5(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[5]),.inputw(inputw12[191:160]),.inputw_index(inputw12_index[39:20]),.counter(`counter),.output_onebank(temp12_result_32[5]));
sparse_mxv sparse12_mxv6(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[6]),.inputw(inputw12[223:192]),.inputw_index(inputw12_index[39:20]),.counter(`counter),.output_onebank(temp12_result_32[6]));
sparse_mxv sparse12_mxv7(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[7]),.inputw(inputw12[255:224]),.inputw_index(inputw12_index[39:20]),.counter(`counter),.output_onebank(temp12_result_32[7]));
sparse_mxv sparse12_mxv8(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[8]),.inputw(inputw12[287:256]),.inputw_index(inputw12_index[59:40]),.counter(`counter),.output_onebank(temp12_result_32[8]));
sparse_mxv sparse12_mxv9(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[9]),.inputw(inputw12[319:288]),.inputw_index(inputw12_index[59:40]),.counter(`counter),.output_onebank(temp12_result_32[9]));
sparse_mxv sparse12_mxv10(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[10]),.inputw(inputw12[351:320]),.inputw_index(inputw12_index[59:40]),.counter(`counter),.output_onebank(temp12_result_32[10]));
sparse_mxv sparse12_mxv11(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[11]),.inputw(inputw12[383:352]),.inputw_index(inputw12_index[59:40]),.counter(`counter),.output_onebank(temp12_result_32[11]));
sparse_mxv sparse12_mxv12(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[12]),.inputw(inputw12[415:384]),.inputw_index(inputw12_index[79:60]),.counter(`counter),.output_onebank(temp12_result_32[12]));
sparse_mxv sparse12_mxv13(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[13]),.inputw(inputw12[447:416]),.inputw_index(inputw12_index[79:60]),.counter(`counter),.output_onebank(temp12_result_32[13]));
sparse_mxv sparse12_mxv14(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[14]),.inputw(inputw12[479:448]),.inputw_index(inputw12_index[79:60]),.counter(`counter),.output_onebank(temp12_result_32[14]));
sparse_mxv sparse12_mxv15(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[15]),.inputw(inputw12[511:480]),.inputw_index(inputw12_index[79:60]),.counter(`counter),.output_onebank(temp12_result_32[15]));
sparse_mxv sparse12_mxv16(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[16]),.inputw(inputw12[543:512]),.inputw_index(inputw12_index[99:80]),.counter(`counter),.output_onebank(temp12_result_32[16]));
sparse_mxv sparse12_mxv17(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[17]),.inputw(inputw12[575:544]),.inputw_index(inputw12_index[99:80]),.counter(`counter),.output_onebank(temp12_result_32[17]));
sparse_mxv sparse12_mxv18(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[18]),.inputw(inputw12[607:576]),.inputw_index(inputw12_index[99:80]),.counter(`counter),.output_onebank(temp12_result_32[18]));
sparse_mxv sparse12_mxv19(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[19]),.inputw(inputw12[639:608]),.inputw_index(inputw12_index[99:80]),.counter(`counter),.output_onebank(temp12_result_32[19]));
sparse_mxv sparse12_mxv20(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[20]),.inputw(inputw12[671:640]),.inputw_index(inputw12_index[119:100]),.counter(`counter),.output_onebank(temp12_result_32[20]));
sparse_mxv sparse12_mxv21(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[21]),.inputw(inputw12[703:672]),.inputw_index(inputw12_index[119:100]),.counter(`counter),.output_onebank(temp12_result_32[21]));
sparse_mxv sparse12_mxv22(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[22]),.inputw(inputw12[735:704]),.inputw_index(inputw12_index[119:100]),.counter(`counter),.output_onebank(temp12_result_32[22]));
sparse_mxv sparse12_mxv23(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[23]),.inputw(inputw12[767:736]),.inputw_index(inputw12_index[119:100]),.counter(`counter),.output_onebank(temp12_result_32[23]));
sparse_mxv sparse12_mxv24(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[24]),.inputw(inputw12[799:768]),.inputw_index(inputw12_index[139:120]),.counter(`counter),.output_onebank(temp12_result_32[24]));
sparse_mxv sparse12_mxv25(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[25]),.inputw(inputw12[831:800]),.inputw_index(inputw12_index[139:120]),.counter(`counter),.output_onebank(temp12_result_32[25]));
sparse_mxv sparse12_mxv26(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[26]),.inputw(inputw12[863:832]),.inputw_index(inputw12_index[139:120]),.counter(`counter),.output_onebank(temp12_result_32[26]));
sparse_mxv sparse12_mxv27(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[27]),.inputw(inputw12[895:864]),.inputw_index(inputw12_index[139:120]),.counter(`counter),.output_onebank(temp12_result_32[27]));
sparse_mxv sparse12_mxv28(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[28]),.inputw(inputw12[927:896]),.inputw_index(inputw12_index[159:140]),.counter(`counter),.output_onebank(temp12_result_32[28]));
sparse_mxv sparse12_mxv29(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[29]),.inputw(inputw12[959:928]),.inputw_index(inputw12_index[159:140]),.counter(`counter),.output_onebank(temp12_result_32[29]));
sparse_mxv sparse12_mxv30(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[30]),.inputw(inputw12[991:960]),.inputw_index(inputw12_index[159:140]),.counter(`counter),.output_onebank(temp12_result_32[30]));
sparse_mxv sparse12_mxv31(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[31]),.inputw(inputw12[1023:992]),.inputw_index(inputw12_index[159:140]),.counter(`counter),.output_onebank(temp12_result_32[31]));
sparse_mxv sparse13_mxv0(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[0]),.inputw(inputw13[31:0]),.inputw_index(inputw13_index[19:0]),.counter(`counter),.output_onebank(temp13_result_32[0]));
sparse_mxv sparse13_mxv1(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[1]),.inputw(inputw13[63:32]),.inputw_index(inputw13_index[19:0]),.counter(`counter),.output_onebank(temp13_result_32[1]));
sparse_mxv sparse13_mxv2(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[2]),.inputw(inputw13[95:64]),.inputw_index(inputw13_index[19:0]),.counter(`counter),.output_onebank(temp13_result_32[2]));
sparse_mxv sparse13_mxv3(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[3]),.inputw(inputw13[127:96]),.inputw_index(inputw13_index[19:0]),.counter(`counter),.output_onebank(temp13_result_32[3]));
sparse_mxv sparse13_mxv4(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[4]),.inputw(inputw13[159:128]),.inputw_index(inputw13_index[39:20]),.counter(`counter),.output_onebank(temp13_result_32[4]));
sparse_mxv sparse13_mxv5(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[5]),.inputw(inputw13[191:160]),.inputw_index(inputw13_index[39:20]),.counter(`counter),.output_onebank(temp13_result_32[5]));
sparse_mxv sparse13_mxv6(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[6]),.inputw(inputw13[223:192]),.inputw_index(inputw13_index[39:20]),.counter(`counter),.output_onebank(temp13_result_32[6]));
sparse_mxv sparse13_mxv7(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[7]),.inputw(inputw13[255:224]),.inputw_index(inputw13_index[39:20]),.counter(`counter),.output_onebank(temp13_result_32[7]));
sparse_mxv sparse13_mxv8(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[8]),.inputw(inputw13[287:256]),.inputw_index(inputw13_index[59:40]),.counter(`counter),.output_onebank(temp13_result_32[8]));
sparse_mxv sparse13_mxv9(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[9]),.inputw(inputw13[319:288]),.inputw_index(inputw13_index[59:40]),.counter(`counter),.output_onebank(temp13_result_32[9]));
sparse_mxv sparse13_mxv10(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[10]),.inputw(inputw13[351:320]),.inputw_index(inputw13_index[59:40]),.counter(`counter),.output_onebank(temp13_result_32[10]));
sparse_mxv sparse13_mxv11(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[11]),.inputw(inputw13[383:352]),.inputw_index(inputw13_index[59:40]),.counter(`counter),.output_onebank(temp13_result_32[11]));
sparse_mxv sparse13_mxv12(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[12]),.inputw(inputw13[415:384]),.inputw_index(inputw13_index[79:60]),.counter(`counter),.output_onebank(temp13_result_32[12]));
sparse_mxv sparse13_mxv13(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[13]),.inputw(inputw13[447:416]),.inputw_index(inputw13_index[79:60]),.counter(`counter),.output_onebank(temp13_result_32[13]));
sparse_mxv sparse13_mxv14(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[14]),.inputw(inputw13[479:448]),.inputw_index(inputw13_index[79:60]),.counter(`counter),.output_onebank(temp13_result_32[14]));
sparse_mxv sparse13_mxv15(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[15]),.inputw(inputw13[511:480]),.inputw_index(inputw13_index[79:60]),.counter(`counter),.output_onebank(temp13_result_32[15]));
sparse_mxv sparse13_mxv16(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[16]),.inputw(inputw13[543:512]),.inputw_index(inputw13_index[99:80]),.counter(`counter),.output_onebank(temp13_result_32[16]));
sparse_mxv sparse13_mxv17(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[17]),.inputw(inputw13[575:544]),.inputw_index(inputw13_index[99:80]),.counter(`counter),.output_onebank(temp13_result_32[17]));
sparse_mxv sparse13_mxv18(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[18]),.inputw(inputw13[607:576]),.inputw_index(inputw13_index[99:80]),.counter(`counter),.output_onebank(temp13_result_32[18]));
sparse_mxv sparse13_mxv19(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[19]),.inputw(inputw13[639:608]),.inputw_index(inputw13_index[99:80]),.counter(`counter),.output_onebank(temp13_result_32[19]));
sparse_mxv sparse13_mxv20(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[20]),.inputw(inputw13[671:640]),.inputw_index(inputw13_index[119:100]),.counter(`counter),.output_onebank(temp13_result_32[20]));
sparse_mxv sparse13_mxv21(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[21]),.inputw(inputw13[703:672]),.inputw_index(inputw13_index[119:100]),.counter(`counter),.output_onebank(temp13_result_32[21]));
sparse_mxv sparse13_mxv22(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[22]),.inputw(inputw13[735:704]),.inputw_index(inputw13_index[119:100]),.counter(`counter),.output_onebank(temp13_result_32[22]));
sparse_mxv sparse13_mxv23(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[23]),.inputw(inputw13[767:736]),.inputw_index(inputw13_index[119:100]),.counter(`counter),.output_onebank(temp13_result_32[23]));
sparse_mxv sparse13_mxv24(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[24]),.inputw(inputw13[799:768]),.inputw_index(inputw13_index[139:120]),.counter(`counter),.output_onebank(temp13_result_32[24]));
sparse_mxv sparse13_mxv25(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[25]),.inputw(inputw13[831:800]),.inputw_index(inputw13_index[139:120]),.counter(`counter),.output_onebank(temp13_result_32[25]));
sparse_mxv sparse13_mxv26(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[26]),.inputw(inputw13[863:832]),.inputw_index(inputw13_index[139:120]),.counter(`counter),.output_onebank(temp13_result_32[26]));
sparse_mxv sparse13_mxv27(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[27]),.inputw(inputw13[895:864]),.inputw_index(inputw13_index[139:120]),.counter(`counter),.output_onebank(temp13_result_32[27]));
sparse_mxv sparse13_mxv28(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[28]),.inputw(inputw13[927:896]),.inputw_index(inputw13_index[159:140]),.counter(`counter),.output_onebank(temp13_result_32[28]));
sparse_mxv sparse13_mxv29(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[29]),.inputw(inputw13[959:928]),.inputw_index(inputw13_index[159:140]),.counter(`counter),.output_onebank(temp13_result_32[29]));
sparse_mxv sparse13_mxv30(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[30]),.inputw(inputw13[991:960]),.inputw_index(inputw13_index[159:140]),.counter(`counter),.output_onebank(temp13_result_32[30]));
sparse_mxv sparse13_mxv31(.clk(clk),.idle(spmvidle3),.rst(rst),.inputx(active_xt[31]),.inputw(inputw13[1023:992]),.inputw_index(inputw13_index[159:140]),.counter(`counter),.output_onebank(temp13_result_32[31]));





always @ (posedge clk) begin // state change 
        if(!rst) begin
            state <= Start ;
            statecount <= 'd0 ;
            spmvidle2 <= 1;
            spmvidle1 <= 1;
            spmvidle <= 1;
            spmvidle3<=1;
        end
        else if (idle) begin
            state <= Start ;
            statecount <= 'd0;
            spmvidle2 <= 1;
            spmvidle1 <= 1;
            spmvidle <= 1;
            spmvidle3<=1;
        end
        else begin
            case(state)
            Start:begin
                state <= Load0;
                statecount <= 'd0;
                spmvidle2 <= spmvidle2;
                spmvidle1 <= spmvidle1;
                spmvidle3 <= spmvidle3;
                spmvidle <= spmvidle ;
            end
            Load0:begin
                state <= Load1;
                statecount <= 'd0;
                spmvidle2 <= spmvidle2;
                spmvidle1 <= spmvidle1;
                spmvidle3 <= spmvidle3;
                spmvidle <= spmvidle ;
            end

            Load1:begin   // latency of Load
                if (statecount <1) begin
                    state <= state;
                    statecount <= statecount + 1;
                    spmvidle2 <= spmvidle2;
                    spmvidle1 <= spmvidle1;
                    spmvidle3 <= spmvidle3;
                    spmvidle <= spmvidle ;
                end 
                else begin
                    state <= Load2;
                    statecount <= statecount + 1;
                    spmvidle2 <= spmvidle2;
                    spmvidle1 <= spmvidle1;
                    spmvidle3 <= spmvidle3;
                    spmvidle <= spmvidle ;
                end
                
            end

            Load2:begin   
                if (statecount <14) begin  //  is Load 16 elements  of active_xt
                    state <= state;
                    statecount <= statecount + 1;
                    spmvidle2 <= spmvidle2;
                    spmvidle1 <= spmvidle1;
                    spmvidle3 <= spmvidle3;
                    spmvidle <= spmvidle ;
                end 
                else begin
                    state <= Load3;
                    statecount <= 'd0;
                    spmvidle2 <= spmvidle2;
                    spmvidle1 <= spmvidle1;
                    spmvidle3 <= spmvidle3;
                    spmvidle <= spmvidle ;
                end
                
            end

            Load3:begin
                state <= Load4;
                statecount <= statecount + 1;
                spmvidle2 <= spmvidle2;
                spmvidle1 <= spmvidle1;
                spmvidle3 <= spmvidle3;
                spmvidle <= spmvidle ;
            end

            Load4:begin
                state <= Wait1;
                statecount <= statecount + 1;
                spmvidle2 <= 1;
                spmvidle1 <= 1;
                spmvidle3 <= 1;
                spmvidle <= 1 ;
            end
            

            Wait1:begin   // the latency time of  sparse_mx
                state <= Wait2;
                statecount <= statecount + 1;
                spmvidle2 <= 0;
                spmvidle1 <= 0;
                spmvidle3 <= 0;
                spmvidle <= 0 ;
            end

            Wait2:begin // the latency time of  sparse_mx
                state <= Wait3;
                statecount <= statecount + 1;
                spmvidle2 <= spmvidle2;
                spmvidle1 <= spmvidle1;
                spmvidle3 <= spmvidle3;
                spmvidle <= spmvidle ;
            end

            Wait3:begin  // the latency time of  sparse_mx
                state <= Wait4;
                statecount <= statecount + 1;
                spmvidle2 <= spmvidle2;
                spmvidle1 <= spmvidle1;
                spmvidle3 <= spmvidle3;
                spmvidle <= spmvidle ;
            end

            Wait4:begin  // the latency time of  sparse_mx
                state <= Wait5;
                statecount <= statecount + 1;
                spmvidle2 <= spmvidle2;
                spmvidle1 <= spmvidle1;
                spmvidle3 <= spmvidle3;
                spmvidle <= spmvidle ;
            end

            Wait5:begin  // the latency time of  sparse_mx
                state <= Wait6;
                statecount <= statecount + 1;
                spmvidle2 <= spmvidle2;
                spmvidle1 <= spmvidle1;
                spmvidle3 <= spmvidle3;
                spmvidle <= spmvidle ;
            end

            Wait6:begin  // the latency time of  sparse_mx
                state <= Wait7;
                statecount <= statecount + 1;
                spmvidle2 <= spmvidle2;
                spmvidle1 <= spmvidle1;
                spmvidle3 <= spmvidle3;
                spmvidle <= spmvidle ;
            end
            
            Wait7:begin  // the latency time of  sparse_mx
                state <= Wait_Add128to64;
                statecount <= statecount + 1;
                spmvidle2 <= spmvidle2;
                spmvidle1 <= spmvidle1;
                spmvidle3 <= spmvidle3;
                spmvidle <= spmvidle ;
            end

            Wait_Add128to64:begin
                state <= Wait_Add128to64_64to32;
                statecount <= statecount + 1;
                spmvidle2 <= spmvidle2;
                spmvidle1 <= spmvidle1;
                spmvidle3 <= spmvidle3;
                spmvidle <= spmvidle ;
            end

            Wait_Add128to64_64to32:begin
                state <= Wait_Add128to64_64to32_32to16;
                statecount <= statecount + 1;
                spmvidle2 <= spmvidle2;
                spmvidle1 <= spmvidle1;
                spmvidle3 <= spmvidle3;
                spmvidle <= spmvidle ;
            end

            Wait_Add128to64_64to32_32to16:begin
                state <= Wait_Add128to64_64to32_32to16_16to8;
                statecount <= statecount + 1;
                spmvidle2 <= spmvidle2;
                spmvidle1 <= spmvidle1;
                spmvidle3 <= spmvidle3;
                spmvidle <= spmvidle ;
            end

            Wait_Add128to64_64to32_32to16_16to8:begin
                state <= Wait_Add128to64_64to32_32to16_16to8_8to4;
                statecount <= statecount + 1;
                spmvidle2 <= spmvidle2;
                spmvidle1 <= spmvidle1;
                spmvidle3 <= spmvidle3;
                spmvidle <= spmvidle ;
            end

            Wait_Add128to64_64to32_32to16_16to8_8to4:begin
                state <= Wait_Add128to64_64to32_32to16_16to8_8to4_4to2;
                statecount <= statecount + 1;
                spmvidle2 <= spmvidle2;
                spmvidle1 <= spmvidle1;
                spmvidle3 <= spmvidle3;
                spmvidle <= spmvidle ;
            end

            Wait_Add128to64_64to32_32to16_16to8_8to4_4to2:begin
                state <= Wait_Add128to64_64to32_32to16_16to8_8to4_4to2_2to1;
                statecount <= statecount + 1;
                spmvidle2 <= spmvidle2;
                spmvidle1 <= spmvidle1;
                spmvidle3 <= spmvidle3;
                spmvidle <= spmvidle ;
            end

            Wait_Add128to64_64to32_32to16_16to8_8to4_4to2_2to1:begin
                spmvidle2 <= spmvidle2;
                spmvidle1 <= spmvidle1;
                spmvidle3 <= spmvidle3;
                spmvidle <= spmvidle ;
                if (statecount < `newcounter) begin // is add 2048 elements 
                    state <= state ;
                    statecount <= statecount + 1;
                end
                else begin
                     state <=Add128to64_64to32_32to16_16to8_8to4_4to2_2to1;
                     statecount <= statecount ;
                end
            end

            Add128to64_64to32_32to16_16to8_8to4_4to2_2to1:begin
                state <= Add64to32_32to16_16to8_8to4_4to2_2to1;
                statecount <= statecount;
                spmvidle2 <= spmvidle2;
                spmvidle1 <= spmvidle1;
                spmvidle3 <= spmvidle3;
                spmvidle <= spmvidle ;
            end

            Add64to32_32to16_16to8_8to4_4to2_2to1:begin
                state <= Add32to16_16to8_8to4_4to2_2to1;
                statecount <= statecount;
                spmvidle2 <= spmvidle2;
                spmvidle1 <= spmvidle1;
                spmvidle3 <= spmvidle3;
                spmvidle <= spmvidle ;
            end

            Add32to16_16to8_8to4_4to2_2to1:begin
                state <= Add16to8_8to4_4to2_2to1;
                statecount <= statecount;
                spmvidle2 <= spmvidle2;
                spmvidle1 <= spmvidle1;
                spmvidle3 <= spmvidle3;
                spmvidle <= spmvidle ;
            end

            Add16to8_8to4_4to2_2to1:begin
                state <= Add8to4_4to2_2to1;
                statecount <= statecount;
                spmvidle2 <= spmvidle2;
                spmvidle1 <= spmvidle1;
                spmvidle3 <= spmvidle3;
                spmvidle <= spmvidle ;
            end

            Add8to4_4to2_2to1:begin
                state <= Add4to2_2to1;
                statecount <= statecount;
                spmvidle2 <= spmvidle2;
                spmvidle1 <= spmvidle1;
                spmvidle3 <= spmvidle3;
                spmvidle <= spmvidle ;
            end

            Add4to2_2to1:begin
                state <= Add2to1;
                statecount <= statecount;
                spmvidle2 <= spmvidle2;
                spmvidle1 <= spmvidle1;
                spmvidle3 <= spmvidle3;
                spmvidle <= spmvidle ;
            end
            Add2to1:begin
                state <= Stop;
                statecount <= statecount;
                spmvidle2 <= spmvidle2;
                spmvidle1 <= spmvidle1;
                spmvidle3 <= spmvidle3;
                spmvidle <= spmvidle ;
            end

            Stop:begin
                state <= state;
                statecount <= statecount;
                spmvidle2 <= spmvidle2;
                spmvidle1 <= spmvidle1;
                spmvidle3 <= spmvidle3;
                spmvidle <= spmvidle ;
            end

            default:begin
                state <= state;
                statecount <= statecount;
                spmvidle2 <= spmvidle2;
                spmvidle1 <= spmvidle1;
                spmvidle3 <= spmvidle3;
                spmvidle <= spmvidle ;
            end

            endcase
        end

end

always @ (posedge clk) begin    // the state machine to assign active_xt reg 
        if(!rst) begin
            active_xt[0] <= active_xt[0];
                active_xt[1] <= active_xt[1];
                active_xt[2] <= active_xt[2];
                active_xt[3] <= active_xt[3];
                active_xt[4] <= active_xt[4];
                active_xt[5] <= active_xt[5];
                active_xt[6] <= active_xt[6];
                active_xt[7] <= active_xt[7];
                active_xt[8] <= active_xt[8];
                active_xt[9] <= active_xt[9];
                active_xt[10] <= active_xt[10];
                active_xt[11] <= active_xt[11];
                active_xt[12] <= active_xt[12];
                active_xt[13] <= active_xt[13];
                active_xt[14] <= active_xt[14];
                active_xt[15] <= active_xt[15];
                active_xt[16] <= active_xt[16];
                active_xt[17] <= active_xt[17];
                active_xt[18] <= active_xt[18];
                active_xt[19] <= active_xt[19];
                active_xt[20] <= active_xt[20];
                active_xt[21] <= active_xt[21];
                active_xt[22] <= active_xt[22];
                active_xt[23] <= active_xt[23];
                active_xt[24] <= active_xt[24];
                active_xt[25] <= active_xt[25];
                active_xt[26] <= active_xt[26];
                active_xt[27] <= active_xt[27];
                active_xt[28] <= active_xt[28];
                active_xt[29] <= active_xt[29];
                active_xt[30] <= active_xt[30];
                active_xt[31] <= active_xt[31];
                
        end
        else if (idle) begin
            active_xt[0] <= active_xt[0];
                active_xt[1] <= active_xt[1];
                active_xt[2] <= active_xt[2];
                active_xt[3] <= active_xt[3];
                active_xt[4] <= active_xt[4];
                active_xt[5] <= active_xt[5];
                active_xt[6] <= active_xt[6];
                active_xt[7] <= active_xt[7];
                active_xt[8] <= active_xt[8];
                active_xt[9] <= active_xt[9];
                active_xt[10] <= active_xt[10];
                active_xt[11] <= active_xt[11];
                active_xt[12] <= active_xt[12];
                active_xt[13] <= active_xt[13];
                active_xt[14] <= active_xt[14];
                active_xt[15] <= active_xt[15];
                active_xt[16] <= active_xt[16];
                active_xt[17] <= active_xt[17];
                active_xt[18] <= active_xt[18];
                active_xt[19] <= active_xt[19];
                active_xt[20] <= active_xt[20];
                active_xt[21] <= active_xt[21];
                active_xt[22] <= active_xt[22];
                active_xt[23] <= active_xt[23];
                active_xt[24] <= active_xt[24];
                active_xt[25] <= active_xt[25];
                
        end
        else begin
            case(state)
            Load2:begin
                if (statecount == 2) begin
                    active_xt[0] <= inputx_output[511:0];
                    active_xt[1] <= inputx_output[1023:512];
                end
                else if (statecount == 3) begin
                    active_xt[2] <= inputx_output[511:0];
                    active_xt[3] <= inputx_output[1023:512];
                end
                else if (statecount == 4) begin
                    active_xt[4] <= inputx_output[511:0];
                    active_xt[5] <= inputx_output[1023:512];
                end
                else if (statecount == 5) begin
                    active_xt[6] <= inputx_output[511:0];
                    active_xt[7] <= inputx_output[1023:512];
                end
                else if (statecount == 6) begin
                    active_xt[8] <= inputx_output[511:0];
                    active_xt[9] <= inputx_output[1023:512];
                end
                else if (statecount == 7) begin
                    active_xt[10] <= inputx_output[511:0];
                    active_xt[11] <= inputx_output[1023:512];
                end
                else if (statecount == 8) begin
                    active_xt[12] <= inputx_output[511:0];
                    active_xt[13] <= inputx_output[1023:512];
                end
                else if (statecount == 9) begin
                    active_xt[14] <= inputx_output[511:0];
                    active_xt[15] <= inputx_output[1023:512];
                end
                else if (statecount == 10) begin
                    active_xt[16] <= inputx_output[511:0];
                    active_xt[17] <= inputx_output[1023:512];
                end
                else if (statecount == 11) begin
                    active_xt[18] <= inputx_output[511:0];
                    active_xt[19] <= inputx_output[1023:512];
                end
                else if (statecount == 12) begin
                    active_xt[20] <= inputx_output[511:0];
                    active_xt[21] <= inputx_output[1023:512];
                end
                else if (statecount == 13) begin
                    active_xt[22] <= inputx_output[511:0];
                    active_xt[23] <= inputx_output[1023:512];
                end
                else if (statecount == 14) begin
                    active_xt[24] <= inputx_output[511:0];
                    active_xt[25] <= inputx_output[1023:512];
                end
                else begin
                    active_xt[0] <= active_xt[0];
                    active_xt[1] <= active_xt[1];
                    active_xt[2] <= active_xt[2];
                    active_xt[3] <= active_xt[3];
                    active_xt[4] <= active_xt[4];
                    active_xt[5] <= active_xt[5];
                    active_xt[6] <= active_xt[6];
                    active_xt[7] <= active_xt[7];
                    active_xt[8] <= active_xt[8];
                    active_xt[9] <= active_xt[9];
                    active_xt[10] <= active_xt[10];
                    active_xt[11] <= active_xt[11];
                    active_xt[12] <= active_xt[12];
                    active_xt[13] <= active_xt[13];
                    active_xt[14] <= active_xt[14];
                    active_xt[15] <= active_xt[15];
                    active_xt[16] <= active_xt[16];
                    active_xt[17] <= active_xt[17];
                    active_xt[18] <= active_xt[18];
                    active_xt[19] <= active_xt[19];
                    active_xt[20] <= active_xt[20];
                    active_xt[21] <= active_xt[21];
                    active_xt[22] <= active_xt[22];
                    active_xt[23] <= active_xt[23];
                    active_xt[24] <= active_xt[24];
                    active_xt[25] <= active_xt[25];
                    
                end
            end
            Load3:begin
                active_xt[26] <= inputx_output[511:0];
                active_xt[27] <= inputx_output[1023:512];
            end
            Load4:begin
                active_xt[28] <= inputx_output[511:0];
                active_xt[29] <= inputx_output[1023:512];
            end
            Wait1:begin
                active_xt[30] <= inputx_output[511:0];
                active_xt[31] <= inputx_output[1023:512];
            end
            default:begin
                active_xt[0] <= active_xt[0];
                active_xt[1] <= active_xt[1];
                active_xt[2] <= active_xt[2];
                active_xt[3] <= active_xt[3];
                active_xt[4] <= active_xt[4];
                active_xt[5] <= active_xt[5];
                active_xt[6] <= active_xt[6];
                active_xt[7] <= active_xt[7];
                active_xt[8] <= active_xt[8];
                active_xt[9] <= active_xt[9];
                active_xt[10] <= active_xt[10];
                active_xt[11] <= active_xt[11];
                active_xt[12] <= active_xt[12];
                active_xt[13] <= active_xt[13];
                active_xt[14] <= active_xt[14];
                active_xt[15] <= active_xt[15];
                active_xt[16] <= active_xt[16];
                active_xt[17] <= active_xt[17];
                active_xt[18] <= active_xt[18];
                active_xt[19] <= active_xt[19];
                active_xt[20] <= active_xt[20];
                active_xt[21] <= active_xt[21];
                active_xt[22] <= active_xt[22];
                active_xt[23] <= active_xt[23];
                active_xt[24] <= active_xt[24];
                active_xt[25] <= active_xt[25];
                active_xt[26] <= active_xt[26];
                active_xt[27] <= active_xt[27];
                active_xt[28] <= active_xt[28];
                active_xt[29] <= active_xt[29];
                active_xt[30] <= active_xt[30];
                active_xt[31] <= active_xt[31];
            end
            endcase
        end
end


always @ (posedge clk) begin    // the state machine to add temp_result_16
        if(!rst) begin
            temp0_result_16[0] <= temp0_result_16[0];
            temp0_result_16[1] <= temp0_result_16[1];
            temp0_result_16[2] <= temp0_result_16[2];
            temp0_result_16[3] <= temp0_result_16[3];
            temp0_result_16[4] <= temp0_result_16[4];
            temp0_result_16[5] <= temp0_result_16[5];
            temp0_result_16[6] <= temp0_result_16[6];
            temp0_result_16[7] <= temp0_result_16[7];
            temp0_result_16[8] <= temp0_result_16[8];
            temp0_result_16[9] <= temp0_result_16[9];
            temp0_result_16[10] <= temp0_result_16[10];
            temp0_result_16[11] <= temp0_result_16[11];
            temp0_result_16[12] <= temp0_result_16[12];
            temp0_result_16[13] <= temp0_result_16[13];
            temp0_result_16[14] <= temp0_result_16[14];
            temp0_result_16[15] <= temp0_result_16[15];
            temp1_result_16[0] <= temp1_result_16[0];
            temp1_result_16[1] <= temp1_result_16[1];
            temp1_result_16[2] <= temp1_result_16[2];
            temp1_result_16[3] <= temp1_result_16[3];
            temp1_result_16[4] <= temp1_result_16[4];
            temp1_result_16[5] <= temp1_result_16[5];
            temp1_result_16[6] <= temp1_result_16[6];
            temp1_result_16[7] <= temp1_result_16[7];
            temp1_result_16[8] <= temp1_result_16[8];
            temp1_result_16[9] <= temp1_result_16[9];
            temp1_result_16[10] <= temp1_result_16[10];
            temp1_result_16[11] <= temp1_result_16[11];
            temp1_result_16[12] <= temp1_result_16[12];
            temp1_result_16[13] <= temp1_result_16[13];
            temp1_result_16[14] <= temp1_result_16[14];
            temp1_result_16[15] <= temp1_result_16[15];

            temp4_result_16[0] <= temp4_result_16[0];
            temp4_result_16[1] <= temp4_result_16[1];
            temp4_result_16[2] <= temp4_result_16[2];
            temp4_result_16[3] <= temp4_result_16[3];
            temp4_result_16[4] <= temp4_result_16[4];
            temp4_result_16[5] <= temp4_result_16[5];
            temp4_result_16[6] <= temp4_result_16[6];
            temp4_result_16[7] <= temp4_result_16[7];
            temp4_result_16[8] <= temp4_result_16[8];
            temp4_result_16[9] <= temp4_result_16[9];
            temp4_result_16[10] <= temp4_result_16[10];
            temp4_result_16[11] <= temp4_result_16[11];
            temp4_result_16[12] <= temp4_result_16[12];
            temp4_result_16[13] <= temp4_result_16[13];
            temp4_result_16[14] <= temp4_result_16[14];
            temp4_result_16[15] <= temp4_result_16[15];
            temp5_result_16[0] <= temp5_result_16[0];
            temp5_result_16[1] <= temp5_result_16[1];
            temp5_result_16[2] <= temp5_result_16[2];
            temp5_result_16[3] <= temp5_result_16[3];
            temp5_result_16[4] <= temp5_result_16[4];
            temp5_result_16[5] <= temp5_result_16[5];
            temp5_result_16[6] <= temp5_result_16[6];
            temp5_result_16[7] <= temp5_result_16[7];
            temp5_result_16[8] <= temp5_result_16[8];
            temp5_result_16[9] <= temp5_result_16[9];
            temp5_result_16[10] <= temp5_result_16[10];
            temp5_result_16[11] <= temp5_result_16[11];
            temp5_result_16[12] <= temp5_result_16[12];
            temp5_result_16[13] <= temp5_result_16[13];
            temp5_result_16[14] <= temp5_result_16[14];
            temp5_result_16[15] <= temp5_result_16[15];

            temp8_result_16[0] <= temp8_result_16[0];
            temp8_result_16[1] <= temp8_result_16[1];
            temp8_result_16[2] <= temp8_result_16[2];
            temp8_result_16[3] <= temp8_result_16[3];
            temp8_result_16[4] <= temp8_result_16[4];
            temp8_result_16[5] <= temp8_result_16[5];
            temp8_result_16[6] <= temp8_result_16[6];
            temp8_result_16[7] <= temp8_result_16[7];
            temp8_result_16[8] <= temp8_result_16[8];
            temp8_result_16[9] <= temp8_result_16[9];
            temp8_result_16[10] <= temp8_result_16[10];
            temp8_result_16[11] <= temp8_result_16[11];
            temp8_result_16[12] <= temp8_result_16[12];
            temp8_result_16[13] <= temp8_result_16[13];
            temp8_result_16[14] <= temp8_result_16[14];
            temp8_result_16[15] <= temp8_result_16[15];
            temp9_result_16[0] <= temp9_result_16[0];
            temp9_result_16[1] <= temp9_result_16[1];
            temp9_result_16[2] <= temp9_result_16[2];
            temp9_result_16[3] <= temp9_result_16[3];
            temp9_result_16[4] <= temp9_result_16[4];
            temp9_result_16[5] <= temp9_result_16[5];
            temp9_result_16[6] <= temp9_result_16[6];
            temp9_result_16[7] <= temp9_result_16[7];
            temp9_result_16[8] <= temp9_result_16[8];
            temp9_result_16[9] <= temp9_result_16[9];
            temp9_result_16[10] <= temp9_result_16[10];
            temp9_result_16[11] <= temp9_result_16[11];
            temp9_result_16[12] <= temp9_result_16[12];
            temp9_result_16[13] <= temp9_result_16[13];
            temp9_result_16[14] <= temp9_result_16[14];
            temp9_result_16[15] <= temp9_result_16[15];

            temp12_result_16[0] <= temp12_result_16[0];
            temp12_result_16[1] <= temp12_result_16[1];
            temp12_result_16[2] <= temp12_result_16[2];
            temp12_result_16[3] <= temp12_result_16[3];
            temp12_result_16[4] <= temp12_result_16[4];
            temp12_result_16[5] <= temp12_result_16[5];
            temp12_result_16[6] <= temp12_result_16[6];
            temp12_result_16[7] <= temp12_result_16[7];
            temp12_result_16[8] <= temp12_result_16[8];
            temp12_result_16[9] <= temp12_result_16[9];
            temp12_result_16[10] <= temp12_result_16[10];
            temp12_result_16[11] <= temp12_result_16[11];
            temp12_result_16[12] <= temp12_result_16[12];
            temp12_result_16[13] <= temp12_result_16[13];
            temp12_result_16[14] <= temp12_result_16[14];
            temp12_result_16[15] <= temp12_result_16[15];
            temp13_result_16[0] <= temp13_result_16[0];
            temp13_result_16[1] <= temp13_result_16[1];
            temp13_result_16[2] <= temp13_result_16[2];
            temp13_result_16[3] <= temp13_result_16[3];
            temp13_result_16[4] <= temp13_result_16[4];
            temp13_result_16[5] <= temp13_result_16[5];
            temp13_result_16[6] <= temp13_result_16[6];
            temp13_result_16[7] <= temp13_result_16[7];
            temp13_result_16[8] <= temp13_result_16[8];
            temp13_result_16[9] <= temp13_result_16[9];
            temp13_result_16[10] <= temp13_result_16[10];
            temp13_result_16[11] <= temp13_result_16[11];
            temp13_result_16[12] <= temp13_result_16[12];
            temp13_result_16[13] <= temp13_result_16[13];
            temp13_result_16[14] <= temp13_result_16[14];
            temp13_result_16[15] <= temp13_result_16[15];

        end
        else if (idle) begin
            temp0_result_16[0] <= temp0_result_16[0];
            temp0_result_16[1] <= temp0_result_16[1];
            temp0_result_16[2] <= temp0_result_16[2];
            temp0_result_16[3] <= temp0_result_16[3];
            temp0_result_16[4] <= temp0_result_16[4];
            temp0_result_16[5] <= temp0_result_16[5];
            temp0_result_16[6] <= temp0_result_16[6];
            temp0_result_16[7] <= temp0_result_16[7];
            temp0_result_16[8] <= temp0_result_16[8];
            temp0_result_16[9] <= temp0_result_16[9];
            temp0_result_16[10] <= temp0_result_16[10];
            temp0_result_16[11] <= temp0_result_16[11];
            temp0_result_16[12] <= temp0_result_16[12];
            temp0_result_16[13] <= temp0_result_16[13];
            temp0_result_16[14] <= temp0_result_16[14];
            temp0_result_16[15] <= temp0_result_16[15];
            temp1_result_16[0] <= temp1_result_16[0];
            temp1_result_16[1] <= temp1_result_16[1];
            temp1_result_16[2] <= temp1_result_16[2];
            temp1_result_16[3] <= temp1_result_16[3];
            temp1_result_16[4] <= temp1_result_16[4];
            temp1_result_16[5] <= temp1_result_16[5];
            temp1_result_16[6] <= temp1_result_16[6];
            temp1_result_16[7] <= temp1_result_16[7];
            temp1_result_16[8] <= temp1_result_16[8];
            temp1_result_16[9] <= temp1_result_16[9];
            temp1_result_16[10] <= temp1_result_16[10];
            temp1_result_16[11] <= temp1_result_16[11];
            temp1_result_16[12] <= temp1_result_16[12];
            temp1_result_16[13] <= temp1_result_16[13];
            temp1_result_16[14] <= temp1_result_16[14];
            temp1_result_16[15] <= temp1_result_16[15];

            temp4_result_16[0] <= temp4_result_16[0];
            temp4_result_16[1] <= temp4_result_16[1];
            temp4_result_16[2] <= temp4_result_16[2];
            temp4_result_16[3] <= temp4_result_16[3];
            temp4_result_16[4] <= temp4_result_16[4];
            temp4_result_16[5] <= temp4_result_16[5];
            temp4_result_16[6] <= temp4_result_16[6];
            temp4_result_16[7] <= temp4_result_16[7];
            temp4_result_16[8] <= temp4_result_16[8];
            temp4_result_16[9] <= temp4_result_16[9];
            temp4_result_16[10] <= temp4_result_16[10];
            temp4_result_16[11] <= temp4_result_16[11];
            temp4_result_16[12] <= temp4_result_16[12];
            temp4_result_16[13] <= temp4_result_16[13];
            temp4_result_16[14] <= temp4_result_16[14];
            temp4_result_16[15] <= temp4_result_16[15];
            temp5_result_16[0] <= temp5_result_16[0];
            temp5_result_16[1] <= temp5_result_16[1];
            temp5_result_16[2] <= temp5_result_16[2];
            temp5_result_16[3] <= temp5_result_16[3];
            temp5_result_16[4] <= temp5_result_16[4];
            temp5_result_16[5] <= temp5_result_16[5];
            temp5_result_16[6] <= temp5_result_16[6];
            temp5_result_16[7] <= temp5_result_16[7];
            temp5_result_16[8] <= temp5_result_16[8];
            temp5_result_16[9] <= temp5_result_16[9];
            temp5_result_16[10] <= temp5_result_16[10];
            temp5_result_16[11] <= temp5_result_16[11];
            temp5_result_16[12] <= temp5_result_16[12];
            temp5_result_16[13] <= temp5_result_16[13];
            temp5_result_16[14] <= temp5_result_16[14];
            temp5_result_16[15] <= temp5_result_16[15];

            temp8_result_16[0] <= temp8_result_16[0];
            temp8_result_16[1] <= temp8_result_16[1];
            temp8_result_16[2] <= temp8_result_16[2];
            temp8_result_16[3] <= temp8_result_16[3];
            temp8_result_16[4] <= temp8_result_16[4];
            temp8_result_16[5] <= temp8_result_16[5];
            temp8_result_16[6] <= temp8_result_16[6];
            temp8_result_16[7] <= temp8_result_16[7];
            temp8_result_16[8] <= temp8_result_16[8];
            temp8_result_16[9] <= temp8_result_16[9];
            temp8_result_16[10] <= temp8_result_16[10];
            temp8_result_16[11] <= temp8_result_16[11];
            temp8_result_16[12] <= temp8_result_16[12];
            temp8_result_16[13] <= temp8_result_16[13];
            temp8_result_16[14] <= temp8_result_16[14];
            temp8_result_16[15] <= temp8_result_16[15];
            temp9_result_16[0] <= temp9_result_16[0];
            temp9_result_16[1] <= temp9_result_16[1];
            temp9_result_16[2] <= temp9_result_16[2];
            temp9_result_16[3] <= temp9_result_16[3];
            temp9_result_16[4] <= temp9_result_16[4];
            temp9_result_16[5] <= temp9_result_16[5];
            temp9_result_16[6] <= temp9_result_16[6];
            temp9_result_16[7] <= temp9_result_16[7];
            temp9_result_16[8] <= temp9_result_16[8];
            temp9_result_16[9] <= temp9_result_16[9];
            temp9_result_16[10] <= temp9_result_16[10];
            temp9_result_16[11] <= temp9_result_16[11];
            temp9_result_16[12] <= temp9_result_16[12];
            temp9_result_16[13] <= temp9_result_16[13];
            temp9_result_16[14] <= temp9_result_16[14];
            temp9_result_16[15] <= temp9_result_16[15];

            temp12_result_16[0] <= temp12_result_16[0];
            temp12_result_16[1] <= temp12_result_16[1];
            temp12_result_16[2] <= temp12_result_16[2];
            temp12_result_16[3] <= temp12_result_16[3];
            temp12_result_16[4] <= temp12_result_16[4];
            temp12_result_16[5] <= temp12_result_16[5];
            temp12_result_16[6] <= temp12_result_16[6];
            temp12_result_16[7] <= temp12_result_16[7];
            temp12_result_16[8] <= temp12_result_16[8];
            temp12_result_16[9] <= temp12_result_16[9];
            temp12_result_16[10] <= temp12_result_16[10];
            temp12_result_16[11] <= temp12_result_16[11];
            temp12_result_16[12] <= temp12_result_16[12];
            temp12_result_16[13] <= temp12_result_16[13];
            temp12_result_16[14] <= temp12_result_16[14];
            temp12_result_16[15] <= temp12_result_16[15];
            temp13_result_16[0] <= temp13_result_16[0];
            temp13_result_16[1] <= temp13_result_16[1];
            temp13_result_16[2] <= temp13_result_16[2];
            temp13_result_16[3] <= temp13_result_16[3];
            temp13_result_16[4] <= temp13_result_16[4];
            temp13_result_16[5] <= temp13_result_16[5];
            temp13_result_16[6] <= temp13_result_16[6];
            temp13_result_16[7] <= temp13_result_16[7];
            temp13_result_16[8] <= temp13_result_16[8];
            temp13_result_16[9] <= temp13_result_16[9];
            temp13_result_16[10] <= temp13_result_16[10];
            temp13_result_16[11] <= temp13_result_16[11];
            temp13_result_16[12] <= temp13_result_16[12];
            temp13_result_16[13] <= temp13_result_16[13];
            temp13_result_16[14] <= temp13_result_16[14];
            temp13_result_16[15] <= temp13_result_16[15];
 
        end
        else begin
            case(state)
            Wait_Add128to64_64to32_32to16:begin
                temp0_result_16[0] <= temp0_result_32[0] + temp0_result_32[1];
                temp0_result_16[1] <= temp0_result_32[2] + temp0_result_32[3];
                temp0_result_16[2] <= temp0_result_32[4] + temp0_result_32[5];
                temp0_result_16[3] <= temp0_result_32[6] + temp0_result_32[7];
                temp0_result_16[4] <= temp0_result_32[8] + temp0_result_32[9];
                temp0_result_16[5] <= temp0_result_32[10] + temp0_result_32[11];
                temp0_result_16[6] <= temp0_result_32[12] + temp0_result_32[13];
                temp0_result_16[7] <= temp0_result_32[14] + temp0_result_32[15];
                temp0_result_16[8] <= temp0_result_32[16] + temp0_result_32[17];
                temp0_result_16[9] <= temp0_result_32[18] + temp0_result_32[19];
                temp0_result_16[10] <= temp0_result_32[20] + temp0_result_32[21];
                temp0_result_16[11] <= temp0_result_32[22] + temp0_result_32[23];
                temp0_result_16[12] <= temp0_result_32[24] + temp0_result_32[25];
                temp0_result_16[13] <= temp0_result_32[26] + temp0_result_32[27];
                temp0_result_16[14] <= temp0_result_32[28] + temp0_result_32[29];
                temp0_result_16[15] <= temp0_result_32[30] + temp0_result_32[31];
                temp1_result_16[0] <= temp1_result_32[0] + temp1_result_32[1];
                temp1_result_16[1] <= temp1_result_32[2] + temp1_result_32[3];
                temp1_result_16[2] <= temp1_result_32[4] + temp1_result_32[5];
                temp1_result_16[3] <= temp1_result_32[6] + temp1_result_32[7];
                temp1_result_16[4] <= temp1_result_32[8] + temp1_result_32[9];
                temp1_result_16[5] <= temp1_result_32[10] + temp1_result_32[11];
                temp1_result_16[6] <= temp1_result_32[12] + temp1_result_32[13];
                temp1_result_16[7] <= temp1_result_32[14] + temp1_result_32[15];
                temp1_result_16[8] <= temp1_result_32[16] + temp1_result_32[17];
                temp1_result_16[9] <= temp1_result_32[18] + temp1_result_32[19];
                temp1_result_16[10] <= temp1_result_32[20] + temp1_result_32[21];
                temp1_result_16[11] <= temp1_result_32[22] + temp1_result_32[23];
                temp1_result_16[12] <= temp1_result_32[24] + temp1_result_32[25];
                temp1_result_16[13] <= temp1_result_32[26] + temp1_result_32[27];
                temp1_result_16[14] <= temp1_result_32[28] + temp1_result_32[29];
                temp1_result_16[15] <= temp1_result_32[30] + temp1_result_32[31];
             
                temp4_result_16[0] <= temp4_result_32[0] + temp4_result_32[1];
                temp4_result_16[1] <= temp4_result_32[2] + temp4_result_32[3];
                temp4_result_16[2] <= temp4_result_32[4] + temp4_result_32[5];
                temp4_result_16[3] <= temp4_result_32[6] + temp4_result_32[7];
                temp4_result_16[4] <= temp4_result_32[8] + temp4_result_32[9];
                temp4_result_16[5] <= temp4_result_32[10] + temp4_result_32[11];
                temp4_result_16[6] <= temp4_result_32[12] + temp4_result_32[13];
                temp4_result_16[7] <= temp4_result_32[14] + temp4_result_32[15];
                temp4_result_16[8] <= temp4_result_32[16] + temp4_result_32[17];
                temp4_result_16[9] <= temp4_result_32[18] + temp4_result_32[19];
                temp4_result_16[10] <= temp4_result_32[20] + temp4_result_32[21];
                temp4_result_16[11] <= temp4_result_32[22] + temp4_result_32[23];
                temp4_result_16[12] <= temp4_result_32[24] + temp4_result_32[25];
                temp4_result_16[13] <= temp4_result_32[26] + temp4_result_32[27];
                temp4_result_16[14] <= temp4_result_32[28] + temp4_result_32[29];
                temp4_result_16[15] <= temp4_result_32[30] + temp4_result_32[31];
                temp5_result_16[0] <= temp5_result_32[0] + temp5_result_32[1];
                temp5_result_16[1] <= temp5_result_32[2] + temp5_result_32[3];
                temp5_result_16[2] <= temp5_result_32[4] + temp5_result_32[5];
                temp5_result_16[3] <= temp5_result_32[6] + temp5_result_32[7];
                temp5_result_16[4] <= temp5_result_32[8] + temp5_result_32[9];
                temp5_result_16[5] <= temp5_result_32[10] + temp5_result_32[11];
                temp5_result_16[6] <= temp5_result_32[12] + temp5_result_32[13];
                temp5_result_16[7] <= temp5_result_32[14] + temp5_result_32[15];
                temp5_result_16[8] <= temp5_result_32[16] + temp5_result_32[17];
                temp5_result_16[9] <= temp5_result_32[18] + temp5_result_32[19];
                temp5_result_16[10] <= temp5_result_32[20] + temp5_result_32[21];
                temp5_result_16[11] <= temp5_result_32[22] + temp5_result_32[23];
                temp5_result_16[12] <= temp5_result_32[24] + temp5_result_32[25];
                temp5_result_16[13] <= temp5_result_32[26] + temp5_result_32[27];
                temp5_result_16[14] <= temp5_result_32[28] + temp5_result_32[29];
                temp5_result_16[15] <= temp5_result_32[30] + temp5_result_32[31];
         
                temp8_result_16[0] <= temp8_result_32[0] + temp8_result_32[1];
                temp8_result_16[1] <= temp8_result_32[2] + temp8_result_32[3];
                temp8_result_16[2] <= temp8_result_32[4] + temp8_result_32[5];
                temp8_result_16[3] <= temp8_result_32[6] + temp8_result_32[7];
                temp8_result_16[4] <= temp8_result_32[8] + temp8_result_32[9];
                temp8_result_16[5] <= temp8_result_32[10] + temp8_result_32[11];
                temp8_result_16[6] <= temp8_result_32[12] + temp8_result_32[13];
                temp8_result_16[7] <= temp8_result_32[14] + temp8_result_32[15];
                temp8_result_16[8] <= temp8_result_32[16] + temp8_result_32[17];
                temp8_result_16[9] <= temp8_result_32[18] + temp8_result_32[19];
                temp8_result_16[10] <= temp8_result_32[20] + temp8_result_32[21];
                temp8_result_16[11] <= temp8_result_32[22] + temp8_result_32[23];
                temp8_result_16[12] <= temp8_result_32[24] + temp8_result_32[25];
                temp8_result_16[13] <= temp8_result_32[26] + temp8_result_32[27];
                temp8_result_16[14] <= temp8_result_32[28] + temp8_result_32[29];
                temp8_result_16[15] <= temp8_result_32[30] + temp8_result_32[31];
                temp9_result_16[0] <= temp9_result_32[0] + temp9_result_32[1];
                temp9_result_16[1] <= temp9_result_32[2] + temp9_result_32[3];
                temp9_result_16[2] <= temp9_result_32[4] + temp9_result_32[5];
                temp9_result_16[3] <= temp9_result_32[6] + temp9_result_32[7];
                temp9_result_16[4] <= temp9_result_32[8] + temp9_result_32[9];
                temp9_result_16[5] <= temp9_result_32[10] + temp9_result_32[11];
                temp9_result_16[6] <= temp9_result_32[12] + temp9_result_32[13];
                temp9_result_16[7] <= temp9_result_32[14] + temp9_result_32[15];
                temp9_result_16[8] <= temp9_result_32[16] + temp9_result_32[17];
                temp9_result_16[9] <= temp9_result_32[18] + temp9_result_32[19];
                temp9_result_16[10] <= temp9_result_32[20] + temp9_result_32[21];
                temp9_result_16[11] <= temp9_result_32[22] + temp9_result_32[23];
                temp9_result_16[12] <= temp9_result_32[24] + temp9_result_32[25];
                temp9_result_16[13] <= temp9_result_32[26] + temp9_result_32[27];
                temp9_result_16[14] <= temp9_result_32[28] + temp9_result_32[29];
                temp9_result_16[15] <= temp9_result_32[30] + temp9_result_32[31];
            
                temp12_result_16[0] <= temp12_result_32[0] + temp12_result_32[1];
                temp12_result_16[1] <= temp12_result_32[2] + temp12_result_32[3];
                temp12_result_16[2] <= temp12_result_32[4] + temp12_result_32[5];
                temp12_result_16[3] <= temp12_result_32[6] + temp12_result_32[7];
                temp12_result_16[4] <= temp12_result_32[8] + temp12_result_32[9];
                temp12_result_16[5] <= temp12_result_32[10] + temp12_result_32[11];
                temp12_result_16[6] <= temp12_result_32[12] + temp12_result_32[13];
                temp12_result_16[7] <= temp12_result_32[14] + temp12_result_32[15];
                temp12_result_16[8] <= temp12_result_32[16] + temp12_result_32[17];
                temp12_result_16[9] <= temp12_result_32[18] + temp12_result_32[19];
                temp12_result_16[10] <= temp12_result_32[20] + temp12_result_32[21];
                temp12_result_16[11] <= temp12_result_32[22] + temp12_result_32[23];
                temp12_result_16[12] <= temp12_result_32[24] + temp12_result_32[25];
                temp12_result_16[13] <= temp12_result_32[26] + temp12_result_32[27];
                temp12_result_16[14] <= temp12_result_32[28] + temp12_result_32[29];
                temp12_result_16[15] <= temp12_result_32[30] + temp12_result_32[31];
                temp13_result_16[0] <= temp13_result_32[0] + temp13_result_32[1];
                temp13_result_16[1] <= temp13_result_32[2] + temp13_result_32[3];
                temp13_result_16[2] <= temp13_result_32[4] + temp13_result_32[5];
                temp13_result_16[3] <= temp13_result_32[6] + temp13_result_32[7];
                temp13_result_16[4] <= temp13_result_32[8] + temp13_result_32[9];
                temp13_result_16[5] <= temp13_result_32[10] + temp13_result_32[11];
                temp13_result_16[6] <= temp13_result_32[12] + temp13_result_32[13];
                temp13_result_16[7] <= temp13_result_32[14] + temp13_result_32[15];
                temp13_result_16[8] <= temp13_result_32[16] + temp13_result_32[17];
                temp13_result_16[9] <= temp13_result_32[18] + temp13_result_32[19];
                temp13_result_16[10] <= temp13_result_32[20] + temp13_result_32[21];
                temp13_result_16[11] <= temp13_result_32[22] + temp13_result_32[23];
                temp13_result_16[12] <= temp13_result_32[24] + temp13_result_32[25];
                temp13_result_16[13] <= temp13_result_32[26] + temp13_result_32[27];
                temp13_result_16[14] <= temp13_result_32[28] + temp13_result_32[29];
                temp13_result_16[15] <= temp13_result_32[30] + temp13_result_32[31];
              
            end
            
            Wait_Add128to64_64to32_32to16_16to8_8to4:begin
                temp0_result_16[0] <= temp0_result_32[0] + temp0_result_32[1];
                temp0_result_16[1] <= temp0_result_32[2] + temp0_result_32[3];
                temp0_result_16[2] <= temp0_result_32[4] + temp0_result_32[5];
                temp0_result_16[3] <= temp0_result_32[6] + temp0_result_32[7];
                temp0_result_16[4] <= temp0_result_32[8] + temp0_result_32[9];
                temp0_result_16[5] <= temp0_result_32[10] + temp0_result_32[11];
                temp0_result_16[6] <= temp0_result_32[12] + temp0_result_32[13];
                temp0_result_16[7] <= temp0_result_32[14] + temp0_result_32[15];
                temp0_result_16[8] <= temp0_result_32[16] + temp0_result_32[17];
                temp0_result_16[9] <= temp0_result_32[18] + temp0_result_32[19];
                temp0_result_16[10] <= temp0_result_32[20] + temp0_result_32[21];
                temp0_result_16[11] <= temp0_result_32[22] + temp0_result_32[23];
                temp0_result_16[12] <= temp0_result_32[24] + temp0_result_32[25];
                temp0_result_16[13] <= temp0_result_32[26] + temp0_result_32[27];
                temp0_result_16[14] <= temp0_result_32[28] + temp0_result_32[29];
                temp0_result_16[15] <= temp0_result_32[30] + temp0_result_32[31];
                temp1_result_16[0] <= temp1_result_32[0] + temp1_result_32[1];
                temp1_result_16[1] <= temp1_result_32[2] + temp1_result_32[3];
                temp1_result_16[2] <= temp1_result_32[4] + temp1_result_32[5];
                temp1_result_16[3] <= temp1_result_32[6] + temp1_result_32[7];
                temp1_result_16[4] <= temp1_result_32[8] + temp1_result_32[9];
                temp1_result_16[5] <= temp1_result_32[10] + temp1_result_32[11];
                temp1_result_16[6] <= temp1_result_32[12] + temp1_result_32[13];
                temp1_result_16[7] <= temp1_result_32[14] + temp1_result_32[15];
                temp1_result_16[8] <= temp1_result_32[16] + temp1_result_32[17];
                temp1_result_16[9] <= temp1_result_32[18] + temp1_result_32[19];
                temp1_result_16[10] <= temp1_result_32[20] + temp1_result_32[21];
                temp1_result_16[11] <= temp1_result_32[22] + temp1_result_32[23];
                temp1_result_16[12] <= temp1_result_32[24] + temp1_result_32[25];
                temp1_result_16[13] <= temp1_result_32[26] + temp1_result_32[27];
                temp1_result_16[14] <= temp1_result_32[28] + temp1_result_32[29];
                temp1_result_16[15] <= temp1_result_32[30] + temp1_result_32[31];
                
                temp4_result_16[0] <= temp4_result_32[0] + temp4_result_32[1];
                temp4_result_16[1] <= temp4_result_32[2] + temp4_result_32[3];
                temp4_result_16[2] <= temp4_result_32[4] + temp4_result_32[5];
                temp4_result_16[3] <= temp4_result_32[6] + temp4_result_32[7];
                temp4_result_16[4] <= temp4_result_32[8] + temp4_result_32[9];
                temp4_result_16[5] <= temp4_result_32[10] + temp4_result_32[11];
                temp4_result_16[6] <= temp4_result_32[12] + temp4_result_32[13];
                temp4_result_16[7] <= temp4_result_32[14] + temp4_result_32[15];
                temp4_result_16[8] <= temp4_result_32[16] + temp4_result_32[17];
                temp4_result_16[9] <= temp4_result_32[18] + temp4_result_32[19];
                temp4_result_16[10] <= temp4_result_32[20] + temp4_result_32[21];
                temp4_result_16[11] <= temp4_result_32[22] + temp4_result_32[23];
                temp4_result_16[12] <= temp4_result_32[24] + temp4_result_32[25];
                temp4_result_16[13] <= temp4_result_32[26] + temp4_result_32[27];
                temp4_result_16[14] <= temp4_result_32[28] + temp4_result_32[29];
                temp4_result_16[15] <= temp4_result_32[30] + temp4_result_32[31];
                temp5_result_16[0] <= temp5_result_32[0] + temp5_result_32[1];
                temp5_result_16[1] <= temp5_result_32[2] + temp5_result_32[3];
                temp5_result_16[2] <= temp5_result_32[4] + temp5_result_32[5];
                temp5_result_16[3] <= temp5_result_32[6] + temp5_result_32[7];
                temp5_result_16[4] <= temp5_result_32[8] + temp5_result_32[9];
                temp5_result_16[5] <= temp5_result_32[10] + temp5_result_32[11];
                temp5_result_16[6] <= temp5_result_32[12] + temp5_result_32[13];
                temp5_result_16[7] <= temp5_result_32[14] + temp5_result_32[15];
                temp5_result_16[8] <= temp5_result_32[16] + temp5_result_32[17];
                temp5_result_16[9] <= temp5_result_32[18] + temp5_result_32[19];
                temp5_result_16[10] <= temp5_result_32[20] + temp5_result_32[21];
                temp5_result_16[11] <= temp5_result_32[22] + temp5_result_32[23];
                temp5_result_16[12] <= temp5_result_32[24] + temp5_result_32[25];
                temp5_result_16[13] <= temp5_result_32[26] + temp5_result_32[27];
                temp5_result_16[14] <= temp5_result_32[28] + temp5_result_32[29];
                temp5_result_16[15] <= temp5_result_32[30] + temp5_result_32[31];
                
                temp8_result_16[0] <= temp8_result_32[0] + temp8_result_32[1];
                temp8_result_16[1] <= temp8_result_32[2] + temp8_result_32[3];
                temp8_result_16[2] <= temp8_result_32[4] + temp8_result_32[5];
                temp8_result_16[3] <= temp8_result_32[6] + temp8_result_32[7];
                temp8_result_16[4] <= temp8_result_32[8] + temp8_result_32[9];
                temp8_result_16[5] <= temp8_result_32[10] + temp8_result_32[11];
                temp8_result_16[6] <= temp8_result_32[12] + temp8_result_32[13];
                temp8_result_16[7] <= temp8_result_32[14] + temp8_result_32[15];
                temp8_result_16[8] <= temp8_result_32[16] + temp8_result_32[17];
                temp8_result_16[9] <= temp8_result_32[18] + temp8_result_32[19];
                temp8_result_16[10] <= temp8_result_32[20] + temp8_result_32[21];
                temp8_result_16[11] <= temp8_result_32[22] + temp8_result_32[23];
                temp8_result_16[12] <= temp8_result_32[24] + temp8_result_32[25];
                temp8_result_16[13] <= temp8_result_32[26] + temp8_result_32[27];
                temp8_result_16[14] <= temp8_result_32[28] + temp8_result_32[29];
                temp8_result_16[15] <= temp8_result_32[30] + temp8_result_32[31];
                temp9_result_16[0] <= temp9_result_32[0] + temp9_result_32[1];
                temp9_result_16[1] <= temp9_result_32[2] + temp9_result_32[3];
                temp9_result_16[2] <= temp9_result_32[4] + temp9_result_32[5];
                temp9_result_16[3] <= temp9_result_32[6] + temp9_result_32[7];
                temp9_result_16[4] <= temp9_result_32[8] + temp9_result_32[9];
                temp9_result_16[5] <= temp9_result_32[10] + temp9_result_32[11];
                temp9_result_16[6] <= temp9_result_32[12] + temp9_result_32[13];
                temp9_result_16[7] <= temp9_result_32[14] + temp9_result_32[15];
                temp9_result_16[8] <= temp9_result_32[16] + temp9_result_32[17];
                temp9_result_16[9] <= temp9_result_32[18] + temp9_result_32[19];
                temp9_result_16[10] <= temp9_result_32[20] + temp9_result_32[21];
                temp9_result_16[11] <= temp9_result_32[22] + temp9_result_32[23];
                temp9_result_16[12] <= temp9_result_32[24] + temp9_result_32[25];
                temp9_result_16[13] <= temp9_result_32[26] + temp9_result_32[27];
                temp9_result_16[14] <= temp9_result_32[28] + temp9_result_32[29];
                temp9_result_16[15] <= temp9_result_32[30] + temp9_result_32[31];
                
                temp12_result_16[0] <= temp12_result_32[0] + temp12_result_32[1];
                temp12_result_16[1] <= temp12_result_32[2] + temp12_result_32[3];
                temp12_result_16[2] <= temp12_result_32[4] + temp12_result_32[5];
                temp12_result_16[3] <= temp12_result_32[6] + temp12_result_32[7];
                temp12_result_16[4] <= temp12_result_32[8] + temp12_result_32[9];
                temp12_result_16[5] <= temp12_result_32[10] + temp12_result_32[11];
                temp12_result_16[6] <= temp12_result_32[12] + temp12_result_32[13];
                temp12_result_16[7] <= temp12_result_32[14] + temp12_result_32[15];
                temp12_result_16[8] <= temp12_result_32[16] + temp12_result_32[17];
                temp12_result_16[9] <= temp12_result_32[18] + temp12_result_32[19];
                temp12_result_16[10] <= temp12_result_32[20] + temp12_result_32[21];
                temp12_result_16[11] <= temp12_result_32[22] + temp12_result_32[23];
                temp12_result_16[12] <= temp12_result_32[24] + temp12_result_32[25];
                temp12_result_16[13] <= temp12_result_32[26] + temp12_result_32[27];
                temp12_result_16[14] <= temp12_result_32[28] + temp12_result_32[29];
                temp12_result_16[15] <= temp12_result_32[30] + temp12_result_32[31];
                temp13_result_16[0] <= temp13_result_32[0] + temp13_result_32[1];
                temp13_result_16[1] <= temp13_result_32[2] + temp13_result_32[3];
                temp13_result_16[2] <= temp13_result_32[4] + temp13_result_32[5];
                temp13_result_16[3] <= temp13_result_32[6] + temp13_result_32[7];
                temp13_result_16[4] <= temp13_result_32[8] + temp13_result_32[9];
                temp13_result_16[5] <= temp13_result_32[10] + temp13_result_32[11];
                temp13_result_16[6] <= temp13_result_32[12] + temp13_result_32[13];
                temp13_result_16[7] <= temp13_result_32[14] + temp13_result_32[15];
                temp13_result_16[8] <= temp13_result_32[16] + temp13_result_32[17];
                temp13_result_16[9] <= temp13_result_32[18] + temp13_result_32[19];
                temp13_result_16[10] <= temp13_result_32[20] + temp13_result_32[21];
                temp13_result_16[11] <= temp13_result_32[22] + temp13_result_32[23];
                temp13_result_16[12] <= temp13_result_32[24] + temp13_result_32[25];
                temp13_result_16[13] <= temp13_result_32[26] + temp13_result_32[27];
                temp13_result_16[14] <= temp13_result_32[28] + temp13_result_32[29];
                temp13_result_16[15] <= temp13_result_32[30] + temp13_result_32[31];
                
            end

            Wait_Add128to64_64to32_32to16_16to8_8to4_4to2:begin
                temp0_result_16[0] <= temp0_result_32[0] + temp0_result_32[1];
                temp0_result_16[1] <= temp0_result_32[2] + temp0_result_32[3];
                temp0_result_16[2] <= temp0_result_32[4] + temp0_result_32[5];
                temp0_result_16[3] <= temp0_result_32[6] + temp0_result_32[7];
                temp0_result_16[4] <= temp0_result_32[8] + temp0_result_32[9];
                temp0_result_16[5] <= temp0_result_32[10] + temp0_result_32[11];
                temp0_result_16[6] <= temp0_result_32[12] + temp0_result_32[13];
                temp0_result_16[7] <= temp0_result_32[14] + temp0_result_32[15];
                temp0_result_16[8] <= temp0_result_32[16] + temp0_result_32[17];
                temp0_result_16[9] <= temp0_result_32[18] + temp0_result_32[19];
                temp0_result_16[10] <= temp0_result_32[20] + temp0_result_32[21];
                temp0_result_16[11] <= temp0_result_32[22] + temp0_result_32[23];
                temp0_result_16[12] <= temp0_result_32[24] + temp0_result_32[25];
                temp0_result_16[13] <= temp0_result_32[26] + temp0_result_32[27];
                temp0_result_16[14] <= temp0_result_32[28] + temp0_result_32[29];
                temp0_result_16[15] <= temp0_result_32[30] + temp0_result_32[31];
                temp1_result_16[0] <= temp1_result_32[0] + temp1_result_32[1];
                temp1_result_16[1] <= temp1_result_32[2] + temp1_result_32[3];
                temp1_result_16[2] <= temp1_result_32[4] + temp1_result_32[5];
                temp1_result_16[3] <= temp1_result_32[6] + temp1_result_32[7];
                temp1_result_16[4] <= temp1_result_32[8] + temp1_result_32[9];
                temp1_result_16[5] <= temp1_result_32[10] + temp1_result_32[11];
                temp1_result_16[6] <= temp1_result_32[12] + temp1_result_32[13];
                temp1_result_16[7] <= temp1_result_32[14] + temp1_result_32[15];
                temp1_result_16[8] <= temp1_result_32[16] + temp1_result_32[17];
                temp1_result_16[9] <= temp1_result_32[18] + temp1_result_32[19];
                temp1_result_16[10] <= temp1_result_32[20] + temp1_result_32[21];
                temp1_result_16[11] <= temp1_result_32[22] + temp1_result_32[23];
                temp1_result_16[12] <= temp1_result_32[24] + temp1_result_32[25];
                temp1_result_16[13] <= temp1_result_32[26] + temp1_result_32[27];
                temp1_result_16[14] <= temp1_result_32[28] + temp1_result_32[29];
                temp1_result_16[15] <= temp1_result_32[30] + temp1_result_32[31];
               
                temp4_result_16[0] <= temp4_result_32[0] + temp4_result_32[1];
                temp4_result_16[1] <= temp4_result_32[2] + temp4_result_32[3];
                temp4_result_16[2] <= temp4_result_32[4] + temp4_result_32[5];
                temp4_result_16[3] <= temp4_result_32[6] + temp4_result_32[7];
                temp4_result_16[4] <= temp4_result_32[8] + temp4_result_32[9];
                temp4_result_16[5] <= temp4_result_32[10] + temp4_result_32[11];
                temp4_result_16[6] <= temp4_result_32[12] + temp4_result_32[13];
                temp4_result_16[7] <= temp4_result_32[14] + temp4_result_32[15];
                temp4_result_16[8] <= temp4_result_32[16] + temp4_result_32[17];
                temp4_result_16[9] <= temp4_result_32[18] + temp4_result_32[19];
                temp4_result_16[10] <= temp4_result_32[20] + temp4_result_32[21];
                temp4_result_16[11] <= temp4_result_32[22] + temp4_result_32[23];
                temp4_result_16[12] <= temp4_result_32[24] + temp4_result_32[25];
                temp4_result_16[13] <= temp4_result_32[26] + temp4_result_32[27];
                temp4_result_16[14] <= temp4_result_32[28] + temp4_result_32[29];
                temp4_result_16[15] <= temp4_result_32[30] + temp4_result_32[31];
                temp5_result_16[0] <= temp5_result_32[0] + temp5_result_32[1];
                temp5_result_16[1] <= temp5_result_32[2] + temp5_result_32[3];
                temp5_result_16[2] <= temp5_result_32[4] + temp5_result_32[5];
                temp5_result_16[3] <= temp5_result_32[6] + temp5_result_32[7];
                temp5_result_16[4] <= temp5_result_32[8] + temp5_result_32[9];
                temp5_result_16[5] <= temp5_result_32[10] + temp5_result_32[11];
                temp5_result_16[6] <= temp5_result_32[12] + temp5_result_32[13];
                temp5_result_16[7] <= temp5_result_32[14] + temp5_result_32[15];
                temp5_result_16[8] <= temp5_result_32[16] + temp5_result_32[17];
                temp5_result_16[9] <= temp5_result_32[18] + temp5_result_32[19];
                temp5_result_16[10] <= temp5_result_32[20] + temp5_result_32[21];
                temp5_result_16[11] <= temp5_result_32[22] + temp5_result_32[23];
                temp5_result_16[12] <= temp5_result_32[24] + temp5_result_32[25];
                temp5_result_16[13] <= temp5_result_32[26] + temp5_result_32[27];
                temp5_result_16[14] <= temp5_result_32[28] + temp5_result_32[29];
                temp5_result_16[15] <= temp5_result_32[30] + temp5_result_32[31];
                
                temp8_result_16[0] <= temp8_result_32[0] + temp8_result_32[1];
                temp8_result_16[1] <= temp8_result_32[2] + temp8_result_32[3];
                temp8_result_16[2] <= temp8_result_32[4] + temp8_result_32[5];
                temp8_result_16[3] <= temp8_result_32[6] + temp8_result_32[7];
                temp8_result_16[4] <= temp8_result_32[8] + temp8_result_32[9];
                temp8_result_16[5] <= temp8_result_32[10] + temp8_result_32[11];
                temp8_result_16[6] <= temp8_result_32[12] + temp8_result_32[13];
                temp8_result_16[7] <= temp8_result_32[14] + temp8_result_32[15];
                temp8_result_16[8] <= temp8_result_32[16] + temp8_result_32[17];
                temp8_result_16[9] <= temp8_result_32[18] + temp8_result_32[19];
                temp8_result_16[10] <= temp8_result_32[20] + temp8_result_32[21];
                temp8_result_16[11] <= temp8_result_32[22] + temp8_result_32[23];
                temp8_result_16[12] <= temp8_result_32[24] + temp8_result_32[25];
                temp8_result_16[13] <= temp8_result_32[26] + temp8_result_32[27];
                temp8_result_16[14] <= temp8_result_32[28] + temp8_result_32[29];
                temp8_result_16[15] <= temp8_result_32[30] + temp8_result_32[31];
                temp9_result_16[0] <= temp9_result_32[0] + temp9_result_32[1];
                temp9_result_16[1] <= temp9_result_32[2] + temp9_result_32[3];
                temp9_result_16[2] <= temp9_result_32[4] + temp9_result_32[5];
                temp9_result_16[3] <= temp9_result_32[6] + temp9_result_32[7];
                temp9_result_16[4] <= temp9_result_32[8] + temp9_result_32[9];
                temp9_result_16[5] <= temp9_result_32[10] + temp9_result_32[11];
                temp9_result_16[6] <= temp9_result_32[12] + temp9_result_32[13];
                temp9_result_16[7] <= temp9_result_32[14] + temp9_result_32[15];
                temp9_result_16[8] <= temp9_result_32[16] + temp9_result_32[17];
                temp9_result_16[9] <= temp9_result_32[18] + temp9_result_32[19];
                temp9_result_16[10] <= temp9_result_32[20] + temp9_result_32[21];
                temp9_result_16[11] <= temp9_result_32[22] + temp9_result_32[23];
                temp9_result_16[12] <= temp9_result_32[24] + temp9_result_32[25];
                temp9_result_16[13] <= temp9_result_32[26] + temp9_result_32[27];
                temp9_result_16[14] <= temp9_result_32[28] + temp9_result_32[29];
                temp9_result_16[15] <= temp9_result_32[30] + temp9_result_32[31];
                
                temp12_result_16[0] <= temp12_result_32[0] + temp12_result_32[1];
                temp12_result_16[1] <= temp12_result_32[2] + temp12_result_32[3];
                temp12_result_16[2] <= temp12_result_32[4] + temp12_result_32[5];
                temp12_result_16[3] <= temp12_result_32[6] + temp12_result_32[7];
                temp12_result_16[4] <= temp12_result_32[8] + temp12_result_32[9];
                temp12_result_16[5] <= temp12_result_32[10] + temp12_result_32[11];
                temp12_result_16[6] <= temp12_result_32[12] + temp12_result_32[13];
                temp12_result_16[7] <= temp12_result_32[14] + temp12_result_32[15];
                temp12_result_16[8] <= temp12_result_32[16] + temp12_result_32[17];
                temp12_result_16[9] <= temp12_result_32[18] + temp12_result_32[19];
                temp12_result_16[10] <= temp12_result_32[20] + temp12_result_32[21];
                temp12_result_16[11] <= temp12_result_32[22] + temp12_result_32[23];
                temp12_result_16[12] <= temp12_result_32[24] + temp12_result_32[25];
                temp12_result_16[13] <= temp12_result_32[26] + temp12_result_32[27];
                temp12_result_16[14] <= temp12_result_32[28] + temp12_result_32[29];
                temp12_result_16[15] <= temp12_result_32[30] + temp12_result_32[31];
                temp13_result_16[0] <= temp13_result_32[0] + temp13_result_32[1];
                temp13_result_16[1] <= temp13_result_32[2] + temp13_result_32[3];
                temp13_result_16[2] <= temp13_result_32[4] + temp13_result_32[5];
                temp13_result_16[3] <= temp13_result_32[6] + temp13_result_32[7];
                temp13_result_16[4] <= temp13_result_32[8] + temp13_result_32[9];
                temp13_result_16[5] <= temp13_result_32[10] + temp13_result_32[11];
                temp13_result_16[6] <= temp13_result_32[12] + temp13_result_32[13];
                temp13_result_16[7] <= temp13_result_32[14] + temp13_result_32[15];
                temp13_result_16[8] <= temp13_result_32[16] + temp13_result_32[17];
                temp13_result_16[9] <= temp13_result_32[18] + temp13_result_32[19];
                temp13_result_16[10] <= temp13_result_32[20] + temp13_result_32[21];
                temp13_result_16[11] <= temp13_result_32[22] + temp13_result_32[23];
                temp13_result_16[12] <= temp13_result_32[24] + temp13_result_32[25];
                temp13_result_16[13] <= temp13_result_32[26] + temp13_result_32[27];
                temp13_result_16[14] <= temp13_result_32[28] + temp13_result_32[29];
                temp13_result_16[15] <= temp13_result_32[30] + temp13_result_32[31];
                
            end

            Wait_Add128to64_64to32_32to16_16to8_8to4_4to2_2to1:begin
                temp0_result_16[0] <= temp0_result_32[0] + temp0_result_32[1];
                temp0_result_16[1] <= temp0_result_32[2] + temp0_result_32[3];
                temp0_result_16[2] <= temp0_result_32[4] + temp0_result_32[5];
                temp0_result_16[3] <= temp0_result_32[6] + temp0_result_32[7];
                temp0_result_16[4] <= temp0_result_32[8] + temp0_result_32[9];
                temp0_result_16[5] <= temp0_result_32[10] + temp0_result_32[11];
                temp0_result_16[6] <= temp0_result_32[12] + temp0_result_32[13];
                temp0_result_16[7] <= temp0_result_32[14] + temp0_result_32[15];
                temp0_result_16[8] <= temp0_result_32[16] + temp0_result_32[17];
                temp0_result_16[9] <= temp0_result_32[18] + temp0_result_32[19];
                temp0_result_16[10] <= temp0_result_32[20] + temp0_result_32[21];
                temp0_result_16[11] <= temp0_result_32[22] + temp0_result_32[23];
                temp0_result_16[12] <= temp0_result_32[24] + temp0_result_32[25];
                temp0_result_16[13] <= temp0_result_32[26] + temp0_result_32[27];
                temp0_result_16[14] <= temp0_result_32[28] + temp0_result_32[29];
                temp0_result_16[15] <= temp0_result_32[30] + temp0_result_32[31];
                temp1_result_16[0] <= temp1_result_32[0] + temp1_result_32[1];
                temp1_result_16[1] <= temp1_result_32[2] + temp1_result_32[3];
                temp1_result_16[2] <= temp1_result_32[4] + temp1_result_32[5];
                temp1_result_16[3] <= temp1_result_32[6] + temp1_result_32[7];
                temp1_result_16[4] <= temp1_result_32[8] + temp1_result_32[9];
                temp1_result_16[5] <= temp1_result_32[10] + temp1_result_32[11];
                temp1_result_16[6] <= temp1_result_32[12] + temp1_result_32[13];
                temp1_result_16[7] <= temp1_result_32[14] + temp1_result_32[15];
                temp1_result_16[8] <= temp1_result_32[16] + temp1_result_32[17];
                temp1_result_16[9] <= temp1_result_32[18] + temp1_result_32[19];
                temp1_result_16[10] <= temp1_result_32[20] + temp1_result_32[21];
                temp1_result_16[11] <= temp1_result_32[22] + temp1_result_32[23];
                temp1_result_16[12] <= temp1_result_32[24] + temp1_result_32[25];
                temp1_result_16[13] <= temp1_result_32[26] + temp1_result_32[27];
                temp1_result_16[14] <= temp1_result_32[28] + temp1_result_32[29];
                temp1_result_16[15] <= temp1_result_32[30] + temp1_result_32[31];
                
                temp4_result_16[0] <= temp4_result_32[0] + temp4_result_32[1];
                temp4_result_16[1] <= temp4_result_32[2] + temp4_result_32[3];
                temp4_result_16[2] <= temp4_result_32[4] + temp4_result_32[5];
                temp4_result_16[3] <= temp4_result_32[6] + temp4_result_32[7];
                temp4_result_16[4] <= temp4_result_32[8] + temp4_result_32[9];
                temp4_result_16[5] <= temp4_result_32[10] + temp4_result_32[11];
                temp4_result_16[6] <= temp4_result_32[12] + temp4_result_32[13];
                temp4_result_16[7] <= temp4_result_32[14] + temp4_result_32[15];
                temp4_result_16[8] <= temp4_result_32[16] + temp4_result_32[17];
                temp4_result_16[9] <= temp4_result_32[18] + temp4_result_32[19];
                temp4_result_16[10] <= temp4_result_32[20] + temp4_result_32[21];
                temp4_result_16[11] <= temp4_result_32[22] + temp4_result_32[23];
                temp4_result_16[12] <= temp4_result_32[24] + temp4_result_32[25];
                temp4_result_16[13] <= temp4_result_32[26] + temp4_result_32[27];
                temp4_result_16[14] <= temp4_result_32[28] + temp4_result_32[29];
                temp4_result_16[15] <= temp4_result_32[30] + temp4_result_32[31];
                temp5_result_16[0] <= temp5_result_32[0] + temp5_result_32[1];
                temp5_result_16[1] <= temp5_result_32[2] + temp5_result_32[3];
                temp5_result_16[2] <= temp5_result_32[4] + temp5_result_32[5];
                temp5_result_16[3] <= temp5_result_32[6] + temp5_result_32[7];
                temp5_result_16[4] <= temp5_result_32[8] + temp5_result_32[9];
                temp5_result_16[5] <= temp5_result_32[10] + temp5_result_32[11];
                temp5_result_16[6] <= temp5_result_32[12] + temp5_result_32[13];
                temp5_result_16[7] <= temp5_result_32[14] + temp5_result_32[15];
                temp5_result_16[8] <= temp5_result_32[16] + temp5_result_32[17];
                temp5_result_16[9] <= temp5_result_32[18] + temp5_result_32[19];
                temp5_result_16[10] <= temp5_result_32[20] + temp5_result_32[21];
                temp5_result_16[11] <= temp5_result_32[22] + temp5_result_32[23];
                temp5_result_16[12] <= temp5_result_32[24] + temp5_result_32[25];
                temp5_result_16[13] <= temp5_result_32[26] + temp5_result_32[27];
                temp5_result_16[14] <= temp5_result_32[28] + temp5_result_32[29];
                temp5_result_16[15] <= temp5_result_32[30] + temp5_result_32[31];
                
                temp8_result_16[0] <= temp8_result_32[0] + temp8_result_32[1];
                temp8_result_16[1] <= temp8_result_32[2] + temp8_result_32[3];
                temp8_result_16[2] <= temp8_result_32[4] + temp8_result_32[5];
                temp8_result_16[3] <= temp8_result_32[6] + temp8_result_32[7];
                temp8_result_16[4] <= temp8_result_32[8] + temp8_result_32[9];
                temp8_result_16[5] <= temp8_result_32[10] + temp8_result_32[11];
                temp8_result_16[6] <= temp8_result_32[12] + temp8_result_32[13];
                temp8_result_16[7] <= temp8_result_32[14] + temp8_result_32[15];
                temp8_result_16[8] <= temp8_result_32[16] + temp8_result_32[17];
                temp8_result_16[9] <= temp8_result_32[18] + temp8_result_32[19];
                temp8_result_16[10] <= temp8_result_32[20] + temp8_result_32[21];
                temp8_result_16[11] <= temp8_result_32[22] + temp8_result_32[23];
                temp8_result_16[12] <= temp8_result_32[24] + temp8_result_32[25];
                temp8_result_16[13] <= temp8_result_32[26] + temp8_result_32[27];
                temp8_result_16[14] <= temp8_result_32[28] + temp8_result_32[29];
                temp8_result_16[15] <= temp8_result_32[30] + temp8_result_32[31];
                temp9_result_16[0] <= temp9_result_32[0] + temp9_result_32[1];
                temp9_result_16[1] <= temp9_result_32[2] + temp9_result_32[3];
                temp9_result_16[2] <= temp9_result_32[4] + temp9_result_32[5];
                temp9_result_16[3] <= temp9_result_32[6] + temp9_result_32[7];
                temp9_result_16[4] <= temp9_result_32[8] + temp9_result_32[9];
                temp9_result_16[5] <= temp9_result_32[10] + temp9_result_32[11];
                temp9_result_16[6] <= temp9_result_32[12] + temp9_result_32[13];
                temp9_result_16[7] <= temp9_result_32[14] + temp9_result_32[15];
                temp9_result_16[8] <= temp9_result_32[16] + temp9_result_32[17];
                temp9_result_16[9] <= temp9_result_32[18] + temp9_result_32[19];
                temp9_result_16[10] <= temp9_result_32[20] + temp9_result_32[21];
                temp9_result_16[11] <= temp9_result_32[22] + temp9_result_32[23];
                temp9_result_16[12] <= temp9_result_32[24] + temp9_result_32[25];
                temp9_result_16[13] <= temp9_result_32[26] + temp9_result_32[27];
                temp9_result_16[14] <= temp9_result_32[28] + temp9_result_32[29];
                temp9_result_16[15] <= temp9_result_32[30] + temp9_result_32[31];
                
                temp12_result_16[0] <= temp12_result_32[0] + temp12_result_32[1];
                temp12_result_16[1] <= temp12_result_32[2] + temp12_result_32[3];
                temp12_result_16[2] <= temp12_result_32[4] + temp12_result_32[5];
                temp12_result_16[3] <= temp12_result_32[6] + temp12_result_32[7];
                temp12_result_16[4] <= temp12_result_32[8] + temp12_result_32[9];
                temp12_result_16[5] <= temp12_result_32[10] + temp12_result_32[11];
                temp12_result_16[6] <= temp12_result_32[12] + temp12_result_32[13];
                temp12_result_16[7] <= temp12_result_32[14] + temp12_result_32[15];
                temp12_result_16[8] <= temp12_result_32[16] + temp12_result_32[17];
                temp12_result_16[9] <= temp12_result_32[18] + temp12_result_32[19];
                temp12_result_16[10] <= temp12_result_32[20] + temp12_result_32[21];
                temp12_result_16[11] <= temp12_result_32[22] + temp12_result_32[23];
                temp12_result_16[12] <= temp12_result_32[24] + temp12_result_32[25];
                temp12_result_16[13] <= temp12_result_32[26] + temp12_result_32[27];
                temp12_result_16[14] <= temp12_result_32[28] + temp12_result_32[29];
                temp12_result_16[15] <= temp12_result_32[30] + temp12_result_32[31];
                temp13_result_16[0] <= temp13_result_32[0] + temp13_result_32[1];
                temp13_result_16[1] <= temp13_result_32[2] + temp13_result_32[3];
                temp13_result_16[2] <= temp13_result_32[4] + temp13_result_32[5];
                temp13_result_16[3] <= temp13_result_32[6] + temp13_result_32[7];
                temp13_result_16[4] <= temp13_result_32[8] + temp13_result_32[9];
                temp13_result_16[5] <= temp13_result_32[10] + temp13_result_32[11];
                temp13_result_16[6] <= temp13_result_32[12] + temp13_result_32[13];
                temp13_result_16[7] <= temp13_result_32[14] + temp13_result_32[15];
                temp13_result_16[8] <= temp13_result_32[16] + temp13_result_32[17];
                temp13_result_16[9] <= temp13_result_32[18] + temp13_result_32[19];
                temp13_result_16[10] <= temp13_result_32[20] + temp13_result_32[21];
                temp13_result_16[11] <= temp13_result_32[22] + temp13_result_32[23];
                temp13_result_16[12] <= temp13_result_32[24] + temp13_result_32[25];
                temp13_result_16[13] <= temp13_result_32[26] + temp13_result_32[27];
                temp13_result_16[14] <= temp13_result_32[28] + temp13_result_32[29];
                temp13_result_16[15] <= temp13_result_32[30] + temp13_result_32[31];
                
            end
            Add128to64_64to32_32to16_16to8_8to4_4to2_2to1:begin
                temp0_result_16[0] <= temp0_result_32[0] + temp0_result_32[1];
                temp0_result_16[1] <= temp0_result_32[2] + temp0_result_32[3];
                temp0_result_16[2] <= temp0_result_32[4] + temp0_result_32[5];
                temp0_result_16[3] <= temp0_result_32[6] + temp0_result_32[7];
                temp0_result_16[4] <= temp0_result_32[8] + temp0_result_32[9];
                temp0_result_16[5] <= temp0_result_32[10] + temp0_result_32[11];
                temp0_result_16[6] <= temp0_result_32[12] + temp0_result_32[13];
                temp0_result_16[7] <= temp0_result_32[14] + temp0_result_32[15];
                temp0_result_16[8] <= temp0_result_32[16] + temp0_result_32[17];
                temp0_result_16[9] <= temp0_result_32[18] + temp0_result_32[19];
                temp0_result_16[10] <= temp0_result_32[20] + temp0_result_32[21];
                temp0_result_16[11] <= temp0_result_32[22] + temp0_result_32[23];
                temp0_result_16[12] <= temp0_result_32[24] + temp0_result_32[25];
                temp0_result_16[13] <= temp0_result_32[26] + temp0_result_32[27];
                temp0_result_16[14] <= temp0_result_32[28] + temp0_result_32[29];
                temp0_result_16[15] <= temp0_result_32[30] + temp0_result_32[31];
                temp1_result_16[0] <= temp1_result_32[0] + temp1_result_32[1];
                temp1_result_16[1] <= temp1_result_32[2] + temp1_result_32[3];
                temp1_result_16[2] <= temp1_result_32[4] + temp1_result_32[5];
                temp1_result_16[3] <= temp1_result_32[6] + temp1_result_32[7];
                temp1_result_16[4] <= temp1_result_32[8] + temp1_result_32[9];
                temp1_result_16[5] <= temp1_result_32[10] + temp1_result_32[11];
                temp1_result_16[6] <= temp1_result_32[12] + temp1_result_32[13];
                temp1_result_16[7] <= temp1_result_32[14] + temp1_result_32[15];
                temp1_result_16[8] <= temp1_result_32[16] + temp1_result_32[17];
                temp1_result_16[9] <= temp1_result_32[18] + temp1_result_32[19];
                temp1_result_16[10] <= temp1_result_32[20] + temp1_result_32[21];
                temp1_result_16[11] <= temp1_result_32[22] + temp1_result_32[23];
                temp1_result_16[12] <= temp1_result_32[24] + temp1_result_32[25];
                temp1_result_16[13] <= temp1_result_32[26] + temp1_result_32[27];
                temp1_result_16[14] <= temp1_result_32[28] + temp1_result_32[29];
                temp1_result_16[15] <= temp1_result_32[30] + temp1_result_32[31];
                
                temp4_result_16[0] <= temp4_result_32[0] + temp4_result_32[1];
                temp4_result_16[1] <= temp4_result_32[2] + temp4_result_32[3];
                temp4_result_16[2] <= temp4_result_32[4] + temp4_result_32[5];
                temp4_result_16[3] <= temp4_result_32[6] + temp4_result_32[7];
                temp4_result_16[4] <= temp4_result_32[8] + temp4_result_32[9];
                temp4_result_16[5] <= temp4_result_32[10] + temp4_result_32[11];
                temp4_result_16[6] <= temp4_result_32[12] + temp4_result_32[13];
                temp4_result_16[7] <= temp4_result_32[14] + temp4_result_32[15];
                temp4_result_16[8] <= temp4_result_32[16] + temp4_result_32[17];
                temp4_result_16[9] <= temp4_result_32[18] + temp4_result_32[19];
                temp4_result_16[10] <= temp4_result_32[20] + temp4_result_32[21];
                temp4_result_16[11] <= temp4_result_32[22] + temp4_result_32[23];
                temp4_result_16[12] <= temp4_result_32[24] + temp4_result_32[25];
                temp4_result_16[13] <= temp4_result_32[26] + temp4_result_32[27];
                temp4_result_16[14] <= temp4_result_32[28] + temp4_result_32[29];
                temp4_result_16[15] <= temp4_result_32[30] + temp4_result_32[31];
                temp5_result_16[0] <= temp5_result_32[0] + temp5_result_32[1];
                temp5_result_16[1] <= temp5_result_32[2] + temp5_result_32[3];
                temp5_result_16[2] <= temp5_result_32[4] + temp5_result_32[5];
                temp5_result_16[3] <= temp5_result_32[6] + temp5_result_32[7];
                temp5_result_16[4] <= temp5_result_32[8] + temp5_result_32[9];
                temp5_result_16[5] <= temp5_result_32[10] + temp5_result_32[11];
                temp5_result_16[6] <= temp5_result_32[12] + temp5_result_32[13];
                temp5_result_16[7] <= temp5_result_32[14] + temp5_result_32[15];
                temp5_result_16[8] <= temp5_result_32[16] + temp5_result_32[17];
                temp5_result_16[9] <= temp5_result_32[18] + temp5_result_32[19];
                temp5_result_16[10] <= temp5_result_32[20] + temp5_result_32[21];
                temp5_result_16[11] <= temp5_result_32[22] + temp5_result_32[23];
                temp5_result_16[12] <= temp5_result_32[24] + temp5_result_32[25];
                temp5_result_16[13] <= temp5_result_32[26] + temp5_result_32[27];
                temp5_result_16[14] <= temp5_result_32[28] + temp5_result_32[29];
                temp5_result_16[15] <= temp5_result_32[30] + temp5_result_32[31];
                
                temp8_result_16[0] <= temp8_result_32[0] + temp8_result_32[1];
                temp8_result_16[1] <= temp8_result_32[2] + temp8_result_32[3];
                temp8_result_16[2] <= temp8_result_32[4] + temp8_result_32[5];
                temp8_result_16[3] <= temp8_result_32[6] + temp8_result_32[7];
                temp8_result_16[4] <= temp8_result_32[8] + temp8_result_32[9];
                temp8_result_16[5] <= temp8_result_32[10] + temp8_result_32[11];
                temp8_result_16[6] <= temp8_result_32[12] + temp8_result_32[13];
                temp8_result_16[7] <= temp8_result_32[14] + temp8_result_32[15];
                temp8_result_16[8] <= temp8_result_32[16] + temp8_result_32[17];
                temp8_result_16[9] <= temp8_result_32[18] + temp8_result_32[19];
                temp8_result_16[10] <= temp8_result_32[20] + temp8_result_32[21];
                temp8_result_16[11] <= temp8_result_32[22] + temp8_result_32[23];
                temp8_result_16[12] <= temp8_result_32[24] + temp8_result_32[25];
                temp8_result_16[13] <= temp8_result_32[26] + temp8_result_32[27];
                temp8_result_16[14] <= temp8_result_32[28] + temp8_result_32[29];
                temp8_result_16[15] <= temp8_result_32[30] + temp8_result_32[31];
                temp9_result_16[0] <= temp9_result_32[0] + temp9_result_32[1];
                temp9_result_16[1] <= temp9_result_32[2] + temp9_result_32[3];
                temp9_result_16[2] <= temp9_result_32[4] + temp9_result_32[5];
                temp9_result_16[3] <= temp9_result_32[6] + temp9_result_32[7];
                temp9_result_16[4] <= temp9_result_32[8] + temp9_result_32[9];
                temp9_result_16[5] <= temp9_result_32[10] + temp9_result_32[11];
                temp9_result_16[6] <= temp9_result_32[12] + temp9_result_32[13];
                temp9_result_16[7] <= temp9_result_32[14] + temp9_result_32[15];
                temp9_result_16[8] <= temp9_result_32[16] + temp9_result_32[17];
                temp9_result_16[9] <= temp9_result_32[18] + temp9_result_32[19];
                temp9_result_16[10] <= temp9_result_32[20] + temp9_result_32[21];
                temp9_result_16[11] <= temp9_result_32[22] + temp9_result_32[23];
                temp9_result_16[12] <= temp9_result_32[24] + temp9_result_32[25];
                temp9_result_16[13] <= temp9_result_32[26] + temp9_result_32[27];
                temp9_result_16[14] <= temp9_result_32[28] + temp9_result_32[29];
                temp9_result_16[15] <= temp9_result_32[30] + temp9_result_32[31];
                
                temp12_result_16[0] <= temp12_result_32[0] + temp12_result_32[1];
                temp12_result_16[1] <= temp12_result_32[2] + temp12_result_32[3];
                temp12_result_16[2] <= temp12_result_32[4] + temp12_result_32[5];
                temp12_result_16[3] <= temp12_result_32[6] + temp12_result_32[7];
                temp12_result_16[4] <= temp12_result_32[8] + temp12_result_32[9];
                temp12_result_16[5] <= temp12_result_32[10] + temp12_result_32[11];
                temp12_result_16[6] <= temp12_result_32[12] + temp12_result_32[13];
                temp12_result_16[7] <= temp12_result_32[14] + temp12_result_32[15];
                temp12_result_16[8] <= temp12_result_32[16] + temp12_result_32[17];
                temp12_result_16[9] <= temp12_result_32[18] + temp12_result_32[19];
                temp12_result_16[10] <= temp12_result_32[20] + temp12_result_32[21];
                temp12_result_16[11] <= temp12_result_32[22] + temp12_result_32[23];
                temp12_result_16[12] <= temp12_result_32[24] + temp12_result_32[25];
                temp12_result_16[13] <= temp12_result_32[26] + temp12_result_32[27];
                temp12_result_16[14] <= temp12_result_32[28] + temp12_result_32[29];
                temp12_result_16[15] <= temp12_result_32[30] + temp12_result_32[31];
                temp13_result_16[0] <= temp13_result_32[0] + temp13_result_32[1];
                temp13_result_16[1] <= temp13_result_32[2] + temp13_result_32[3];
                temp13_result_16[2] <= temp13_result_32[4] + temp13_result_32[5];
                temp13_result_16[3] <= temp13_result_32[6] + temp13_result_32[7];
                temp13_result_16[4] <= temp13_result_32[8] + temp13_result_32[9];
                temp13_result_16[5] <= temp13_result_32[10] + temp13_result_32[11];
                temp13_result_16[6] <= temp13_result_32[12] + temp13_result_32[13];
                temp13_result_16[7] <= temp13_result_32[14] + temp13_result_32[15];
                temp13_result_16[8] <= temp13_result_32[16] + temp13_result_32[17];
                temp13_result_16[9] <= temp13_result_32[18] + temp13_result_32[19];
                temp13_result_16[10] <= temp13_result_32[20] + temp13_result_32[21];
                temp13_result_16[11] <= temp13_result_32[22] + temp13_result_32[23];
                temp13_result_16[12] <= temp13_result_32[24] + temp13_result_32[25];
                temp13_result_16[13] <= temp13_result_32[26] + temp13_result_32[27];
                temp13_result_16[14] <= temp13_result_32[28] + temp13_result_32[29];
                temp13_result_16[15] <= temp13_result_32[30] + temp13_result_32[31];
                
            end
            Add64to32_32to16_16to8_8to4_4to2_2to1:begin
                temp0_result_16[0] <= temp0_result_32[0] + temp0_result_32[1];
                temp0_result_16[1] <= temp0_result_32[2] + temp0_result_32[3];
                temp0_result_16[2] <= temp0_result_32[4] + temp0_result_32[5];
                temp0_result_16[3] <= temp0_result_32[6] + temp0_result_32[7];
                temp0_result_16[4] <= temp0_result_32[8] + temp0_result_32[9];
                temp0_result_16[5] <= temp0_result_32[10] + temp0_result_32[11];
                temp0_result_16[6] <= temp0_result_32[12] + temp0_result_32[13];
                temp0_result_16[7] <= temp0_result_32[14] + temp0_result_32[15];
                temp0_result_16[8] <= temp0_result_32[16] + temp0_result_32[17];
                temp0_result_16[9] <= temp0_result_32[18] + temp0_result_32[19];
                temp0_result_16[10] <= temp0_result_32[20] + temp0_result_32[21];
                temp0_result_16[11] <= temp0_result_32[22] + temp0_result_32[23];
                temp0_result_16[12] <= temp0_result_32[24] + temp0_result_32[25];
                temp0_result_16[13] <= temp0_result_32[26] + temp0_result_32[27];
                temp0_result_16[14] <= temp0_result_32[28] + temp0_result_32[29];
                temp0_result_16[15] <= temp0_result_32[30] + temp0_result_32[31];
                temp1_result_16[0] <= temp1_result_32[0] + temp1_result_32[1];
                temp1_result_16[1] <= temp1_result_32[2] + temp1_result_32[3];
                temp1_result_16[2] <= temp1_result_32[4] + temp1_result_32[5];
                temp1_result_16[3] <= temp1_result_32[6] + temp1_result_32[7];
                temp1_result_16[4] <= temp1_result_32[8] + temp1_result_32[9];
                temp1_result_16[5] <= temp1_result_32[10] + temp1_result_32[11];
                temp1_result_16[6] <= temp1_result_32[12] + temp1_result_32[13];
                temp1_result_16[7] <= temp1_result_32[14] + temp1_result_32[15];
                temp1_result_16[8] <= temp1_result_32[16] + temp1_result_32[17];
                temp1_result_16[9] <= temp1_result_32[18] + temp1_result_32[19];
                temp1_result_16[10] <= temp1_result_32[20] + temp1_result_32[21];
                temp1_result_16[11] <= temp1_result_32[22] + temp1_result_32[23];
                temp1_result_16[12] <= temp1_result_32[24] + temp1_result_32[25];
                temp1_result_16[13] <= temp1_result_32[26] + temp1_result_32[27];
                temp1_result_16[14] <= temp1_result_32[28] + temp1_result_32[29];
                temp1_result_16[15] <= temp1_result_32[30] + temp1_result_32[31];
                
               
                temp4_result_16[0] <= temp4_result_32[0] + temp4_result_32[1];
                temp4_result_16[1] <= temp4_result_32[2] + temp4_result_32[3];
                temp4_result_16[2] <= temp4_result_32[4] + temp4_result_32[5];
                temp4_result_16[3] <= temp4_result_32[6] + temp4_result_32[7];
                temp4_result_16[4] <= temp4_result_32[8] + temp4_result_32[9];
                temp4_result_16[5] <= temp4_result_32[10] + temp4_result_32[11];
                temp4_result_16[6] <= temp4_result_32[12] + temp4_result_32[13];
                temp4_result_16[7] <= temp4_result_32[14] + temp4_result_32[15];
                temp4_result_16[8] <= temp4_result_32[16] + temp4_result_32[17];
                temp4_result_16[9] <= temp4_result_32[18] + temp4_result_32[19];
                temp4_result_16[10] <= temp4_result_32[20] + temp4_result_32[21];
                temp4_result_16[11] <= temp4_result_32[22] + temp4_result_32[23];
                temp4_result_16[12] <= temp4_result_32[24] + temp4_result_32[25];
                temp4_result_16[13] <= temp4_result_32[26] + temp4_result_32[27];
                temp4_result_16[14] <= temp4_result_32[28] + temp4_result_32[29];
                temp4_result_16[15] <= temp4_result_32[30] + temp4_result_32[31];
                temp5_result_16[0] <= temp5_result_32[0] + temp5_result_32[1];
                temp5_result_16[1] <= temp5_result_32[2] + temp5_result_32[3];
                temp5_result_16[2] <= temp5_result_32[4] + temp5_result_32[5];
                temp5_result_16[3] <= temp5_result_32[6] + temp5_result_32[7];
                temp5_result_16[4] <= temp5_result_32[8] + temp5_result_32[9];
                temp5_result_16[5] <= temp5_result_32[10] + temp5_result_32[11];
                temp5_result_16[6] <= temp5_result_32[12] + temp5_result_32[13];
                temp5_result_16[7] <= temp5_result_32[14] + temp5_result_32[15];
                temp5_result_16[8] <= temp5_result_32[16] + temp5_result_32[17];
                temp5_result_16[9] <= temp5_result_32[18] + temp5_result_32[19];
                temp5_result_16[10] <= temp5_result_32[20] + temp5_result_32[21];
                temp5_result_16[11] <= temp5_result_32[22] + temp5_result_32[23];
                temp5_result_16[12] <= temp5_result_32[24] + temp5_result_32[25];
                temp5_result_16[13] <= temp5_result_32[26] + temp5_result_32[27];
                temp5_result_16[14] <= temp5_result_32[28] + temp5_result_32[29];
                temp5_result_16[15] <= temp5_result_32[30] + temp5_result_32[31];
               
                temp8_result_16[0] <= temp8_result_32[0] + temp8_result_32[1];
                temp8_result_16[1] <= temp8_result_32[2] + temp8_result_32[3];
                temp8_result_16[2] <= temp8_result_32[4] + temp8_result_32[5];
                temp8_result_16[3] <= temp8_result_32[6] + temp8_result_32[7];
                temp8_result_16[4] <= temp8_result_32[8] + temp8_result_32[9];
                temp8_result_16[5] <= temp8_result_32[10] + temp8_result_32[11];
                temp8_result_16[6] <= temp8_result_32[12] + temp8_result_32[13];
                temp8_result_16[7] <= temp8_result_32[14] + temp8_result_32[15];
                temp8_result_16[8] <= temp8_result_32[16] + temp8_result_32[17];
                temp8_result_16[9] <= temp8_result_32[18] + temp8_result_32[19];
                temp8_result_16[10] <= temp8_result_32[20] + temp8_result_32[21];
                temp8_result_16[11] <= temp8_result_32[22] + temp8_result_32[23];
                temp8_result_16[12] <= temp8_result_32[24] + temp8_result_32[25];
                temp8_result_16[13] <= temp8_result_32[26] + temp8_result_32[27];
                temp8_result_16[14] <= temp8_result_32[28] + temp8_result_32[29];
                temp8_result_16[15] <= temp8_result_32[30] + temp8_result_32[31];
                temp9_result_16[0] <= temp9_result_32[0] + temp9_result_32[1];
                temp9_result_16[1] <= temp9_result_32[2] + temp9_result_32[3];
                temp9_result_16[2] <= temp9_result_32[4] + temp9_result_32[5];
                temp9_result_16[3] <= temp9_result_32[6] + temp9_result_32[7];
                temp9_result_16[4] <= temp9_result_32[8] + temp9_result_32[9];
                temp9_result_16[5] <= temp9_result_32[10] + temp9_result_32[11];
                temp9_result_16[6] <= temp9_result_32[12] + temp9_result_32[13];
                temp9_result_16[7] <= temp9_result_32[14] + temp9_result_32[15];
                temp9_result_16[8] <= temp9_result_32[16] + temp9_result_32[17];
                temp9_result_16[9] <= temp9_result_32[18] + temp9_result_32[19];
                temp9_result_16[10] <= temp9_result_32[20] + temp9_result_32[21];
                temp9_result_16[11] <= temp9_result_32[22] + temp9_result_32[23];
                temp9_result_16[12] <= temp9_result_32[24] + temp9_result_32[25];
                temp9_result_16[13] <= temp9_result_32[26] + temp9_result_32[27];
                temp9_result_16[14] <= temp9_result_32[28] + temp9_result_32[29];
                temp9_result_16[15] <= temp9_result_32[30] + temp9_result_32[31];
                
                temp12_result_16[0] <= temp12_result_32[0] + temp12_result_32[1];
                temp12_result_16[1] <= temp12_result_32[2] + temp12_result_32[3];
                temp12_result_16[2] <= temp12_result_32[4] + temp12_result_32[5];
                temp12_result_16[3] <= temp12_result_32[6] + temp12_result_32[7];
                temp12_result_16[4] <= temp12_result_32[8] + temp12_result_32[9];
                temp12_result_16[5] <= temp12_result_32[10] + temp12_result_32[11];
                temp12_result_16[6] <= temp12_result_32[12] + temp12_result_32[13];
                temp12_result_16[7] <= temp12_result_32[14] + temp12_result_32[15];
                temp12_result_16[8] <= temp12_result_32[16] + temp12_result_32[17];
                temp12_result_16[9] <= temp12_result_32[18] + temp12_result_32[19];
                temp12_result_16[10] <= temp12_result_32[20] + temp12_result_32[21];
                temp12_result_16[11] <= temp12_result_32[22] + temp12_result_32[23];
                temp12_result_16[12] <= temp12_result_32[24] + temp12_result_32[25];
                temp12_result_16[13] <= temp12_result_32[26] + temp12_result_32[27];
                temp12_result_16[14] <= temp12_result_32[28] + temp12_result_32[29];
                temp12_result_16[15] <= temp12_result_32[30] + temp12_result_32[31];
                temp13_result_16[0] <= temp13_result_32[0] + temp13_result_32[1];
                temp13_result_16[1] <= temp13_result_32[2] + temp13_result_32[3];
                temp13_result_16[2] <= temp13_result_32[4] + temp13_result_32[5];
                temp13_result_16[3] <= temp13_result_32[6] + temp13_result_32[7];
                temp13_result_16[4] <= temp13_result_32[8] + temp13_result_32[9];
                temp13_result_16[5] <= temp13_result_32[10] + temp13_result_32[11];
                temp13_result_16[6] <= temp13_result_32[12] + temp13_result_32[13];
                temp13_result_16[7] <= temp13_result_32[14] + temp13_result_32[15];
                temp13_result_16[8] <= temp13_result_32[16] + temp13_result_32[17];
                temp13_result_16[9] <= temp13_result_32[18] + temp13_result_32[19];
                temp13_result_16[10] <= temp13_result_32[20] + temp13_result_32[21];
                temp13_result_16[11] <= temp13_result_32[22] + temp13_result_32[23];
                temp13_result_16[12] <= temp13_result_32[24] + temp13_result_32[25];
                temp13_result_16[13] <= temp13_result_32[26] + temp13_result_32[27];
                temp13_result_16[14] <= temp13_result_32[28] + temp13_result_32[29];
                temp13_result_16[15] <= temp13_result_32[30] + temp13_result_32[31];
                
            end
            Add32to16_16to8_8to4_4to2_2to1:begin
                temp0_result_16[0] <= temp0_result_32[0] + temp0_result_32[1];
                temp0_result_16[1] <= temp0_result_32[2] + temp0_result_32[3];
                temp0_result_16[2] <= temp0_result_32[4] + temp0_result_32[5];
                temp0_result_16[3] <= temp0_result_32[6] + temp0_result_32[7];
                temp0_result_16[4] <= temp0_result_32[8] + temp0_result_32[9];
                temp0_result_16[5] <= temp0_result_32[10] + temp0_result_32[11];
                temp0_result_16[6] <= temp0_result_32[12] + temp0_result_32[13];
                temp0_result_16[7] <= temp0_result_32[14] + temp0_result_32[15];
                temp0_result_16[8] <= temp0_result_32[16] + temp0_result_32[17];
                temp0_result_16[9] <= temp0_result_32[18] + temp0_result_32[19];
                temp0_result_16[10] <= temp0_result_32[20] + temp0_result_32[21];
                temp0_result_16[11] <= temp0_result_32[22] + temp0_result_32[23];
                temp0_result_16[12] <= temp0_result_32[24] + temp0_result_32[25];
                temp0_result_16[13] <= temp0_result_32[26] + temp0_result_32[27];
                temp0_result_16[14] <= temp0_result_32[28] + temp0_result_32[29];
                temp0_result_16[15] <= temp0_result_32[30] + temp0_result_32[31];
                temp1_result_16[0] <= temp1_result_32[0] + temp1_result_32[1];
                temp1_result_16[1] <= temp1_result_32[2] + temp1_result_32[3];
                temp1_result_16[2] <= temp1_result_32[4] + temp1_result_32[5];
                temp1_result_16[3] <= temp1_result_32[6] + temp1_result_32[7];
                temp1_result_16[4] <= temp1_result_32[8] + temp1_result_32[9];
                temp1_result_16[5] <= temp1_result_32[10] + temp1_result_32[11];
                temp1_result_16[6] <= temp1_result_32[12] + temp1_result_32[13];
                temp1_result_16[7] <= temp1_result_32[14] + temp1_result_32[15];
                temp1_result_16[8] <= temp1_result_32[16] + temp1_result_32[17];
                temp1_result_16[9] <= temp1_result_32[18] + temp1_result_32[19];
                temp1_result_16[10] <= temp1_result_32[20] + temp1_result_32[21];
                temp1_result_16[11] <= temp1_result_32[22] + temp1_result_32[23];
                temp1_result_16[12] <= temp1_result_32[24] + temp1_result_32[25];
                temp1_result_16[13] <= temp1_result_32[26] + temp1_result_32[27];
                temp1_result_16[14] <= temp1_result_32[28] + temp1_result_32[29];
                temp1_result_16[15] <= temp1_result_32[30] + temp1_result_32[31];
                
               
                temp4_result_16[0] <= temp4_result_32[0] + temp4_result_32[1];
                temp4_result_16[1] <= temp4_result_32[2] + temp4_result_32[3];
                temp4_result_16[2] <= temp4_result_32[4] + temp4_result_32[5];
                temp4_result_16[3] <= temp4_result_32[6] + temp4_result_32[7];
                temp4_result_16[4] <= temp4_result_32[8] + temp4_result_32[9];
                temp4_result_16[5] <= temp4_result_32[10] + temp4_result_32[11];
                temp4_result_16[6] <= temp4_result_32[12] + temp4_result_32[13];
                temp4_result_16[7] <= temp4_result_32[14] + temp4_result_32[15];
                temp4_result_16[8] <= temp4_result_32[16] + temp4_result_32[17];
                temp4_result_16[9] <= temp4_result_32[18] + temp4_result_32[19];
                temp4_result_16[10] <= temp4_result_32[20] + temp4_result_32[21];
                temp4_result_16[11] <= temp4_result_32[22] + temp4_result_32[23];
                temp4_result_16[12] <= temp4_result_32[24] + temp4_result_32[25];
                temp4_result_16[13] <= temp4_result_32[26] + temp4_result_32[27];
                temp4_result_16[14] <= temp4_result_32[28] + temp4_result_32[29];
                temp4_result_16[15] <= temp4_result_32[30] + temp4_result_32[31];
                temp5_result_16[0] <= temp5_result_32[0] + temp5_result_32[1];
                temp5_result_16[1] <= temp5_result_32[2] + temp5_result_32[3];
                temp5_result_16[2] <= temp5_result_32[4] + temp5_result_32[5];
                temp5_result_16[3] <= temp5_result_32[6] + temp5_result_32[7];
                temp5_result_16[4] <= temp5_result_32[8] + temp5_result_32[9];
                temp5_result_16[5] <= temp5_result_32[10] + temp5_result_32[11];
                temp5_result_16[6] <= temp5_result_32[12] + temp5_result_32[13];
                temp5_result_16[7] <= temp5_result_32[14] + temp5_result_32[15];
                temp5_result_16[8] <= temp5_result_32[16] + temp5_result_32[17];
                temp5_result_16[9] <= temp5_result_32[18] + temp5_result_32[19];
                temp5_result_16[10] <= temp5_result_32[20] + temp5_result_32[21];
                temp5_result_16[11] <= temp5_result_32[22] + temp5_result_32[23];
                temp5_result_16[12] <= temp5_result_32[24] + temp5_result_32[25];
                temp5_result_16[13] <= temp5_result_32[26] + temp5_result_32[27];
                temp5_result_16[14] <= temp5_result_32[28] + temp5_result_32[29];
                temp5_result_16[15] <= temp5_result_32[30] + temp5_result_32[31];
               
                temp8_result_16[0] <= temp8_result_32[0] + temp8_result_32[1];
                temp8_result_16[1] <= temp8_result_32[2] + temp8_result_32[3];
                temp8_result_16[2] <= temp8_result_32[4] + temp8_result_32[5];
                temp8_result_16[3] <= temp8_result_32[6] + temp8_result_32[7];
                temp8_result_16[4] <= temp8_result_32[8] + temp8_result_32[9];
                temp8_result_16[5] <= temp8_result_32[10] + temp8_result_32[11];
                temp8_result_16[6] <= temp8_result_32[12] + temp8_result_32[13];
                temp8_result_16[7] <= temp8_result_32[14] + temp8_result_32[15];
                temp8_result_16[8] <= temp8_result_32[16] + temp8_result_32[17];
                temp8_result_16[9] <= temp8_result_32[18] + temp8_result_32[19];
                temp8_result_16[10] <= temp8_result_32[20] + temp8_result_32[21];
                temp8_result_16[11] <= temp8_result_32[22] + temp8_result_32[23];
                temp8_result_16[12] <= temp8_result_32[24] + temp8_result_32[25];
                temp8_result_16[13] <= temp8_result_32[26] + temp8_result_32[27];
                temp8_result_16[14] <= temp8_result_32[28] + temp8_result_32[29];
                temp8_result_16[15] <= temp8_result_32[30] + temp8_result_32[31];
                temp9_result_16[0] <= temp9_result_32[0] + temp9_result_32[1];
                temp9_result_16[1] <= temp9_result_32[2] + temp9_result_32[3];
                temp9_result_16[2] <= temp9_result_32[4] + temp9_result_32[5];
                temp9_result_16[3] <= temp9_result_32[6] + temp9_result_32[7];
                temp9_result_16[4] <= temp9_result_32[8] + temp9_result_32[9];
                temp9_result_16[5] <= temp9_result_32[10] + temp9_result_32[11];
                temp9_result_16[6] <= temp9_result_32[12] + temp9_result_32[13];
                temp9_result_16[7] <= temp9_result_32[14] + temp9_result_32[15];
                temp9_result_16[8] <= temp9_result_32[16] + temp9_result_32[17];
                temp9_result_16[9] <= temp9_result_32[18] + temp9_result_32[19];
                temp9_result_16[10] <= temp9_result_32[20] + temp9_result_32[21];
                temp9_result_16[11] <= temp9_result_32[22] + temp9_result_32[23];
                temp9_result_16[12] <= temp9_result_32[24] + temp9_result_32[25];
                temp9_result_16[13] <= temp9_result_32[26] + temp9_result_32[27];
                temp9_result_16[14] <= temp9_result_32[28] + temp9_result_32[29];
                temp9_result_16[15] <= temp9_result_32[30] + temp9_result_32[31];
                
                temp12_result_16[0] <= temp12_result_32[0] + temp12_result_32[1];
                temp12_result_16[1] <= temp12_result_32[2] + temp12_result_32[3];
                temp12_result_16[2] <= temp12_result_32[4] + temp12_result_32[5];
                temp12_result_16[3] <= temp12_result_32[6] + temp12_result_32[7];
                temp12_result_16[4] <= temp12_result_32[8] + temp12_result_32[9];
                temp12_result_16[5] <= temp12_result_32[10] + temp12_result_32[11];
                temp12_result_16[6] <= temp12_result_32[12] + temp12_result_32[13];
                temp12_result_16[7] <= temp12_result_32[14] + temp12_result_32[15];
                temp12_result_16[8] <= temp12_result_32[16] + temp12_result_32[17];
                temp12_result_16[9] <= temp12_result_32[18] + temp12_result_32[19];
                temp12_result_16[10] <= temp12_result_32[20] + temp12_result_32[21];
                temp12_result_16[11] <= temp12_result_32[22] + temp12_result_32[23];
                temp12_result_16[12] <= temp12_result_32[24] + temp12_result_32[25];
                temp12_result_16[13] <= temp12_result_32[26] + temp12_result_32[27];
                temp12_result_16[14] <= temp12_result_32[28] + temp12_result_32[29];
                temp12_result_16[15] <= temp12_result_32[30] + temp12_result_32[31];
                temp13_result_16[0] <= temp13_result_32[0] + temp13_result_32[1];
                temp13_result_16[1] <= temp13_result_32[2] + temp13_result_32[3];
                temp13_result_16[2] <= temp13_result_32[4] + temp13_result_32[5];
                temp13_result_16[3] <= temp13_result_32[6] + temp13_result_32[7];
                temp13_result_16[4] <= temp13_result_32[8] + temp13_result_32[9];
                temp13_result_16[5] <= temp13_result_32[10] + temp13_result_32[11];
                temp13_result_16[6] <= temp13_result_32[12] + temp13_result_32[13];
                temp13_result_16[7] <= temp13_result_32[14] + temp13_result_32[15];
                temp13_result_16[8] <= temp13_result_32[16] + temp13_result_32[17];
                temp13_result_16[9] <= temp13_result_32[18] + temp13_result_32[19];
                temp13_result_16[10] <= temp13_result_32[20] + temp13_result_32[21];
                temp13_result_16[11] <= temp13_result_32[22] + temp13_result_32[23];
                temp13_result_16[12] <= temp13_result_32[24] + temp13_result_32[25];
                temp13_result_16[13] <= temp13_result_32[26] + temp13_result_32[27];
                temp13_result_16[14] <= temp13_result_32[28] + temp13_result_32[29];
                temp13_result_16[15] <= temp13_result_32[30] + temp13_result_32[31];
            end
            default:begin
                temp0_result_16[0] <= temp0_result_16[0];
            temp0_result_16[1] <= temp0_result_16[1];
            temp0_result_16[2] <= temp0_result_16[2];
            temp0_result_16[3] <= temp0_result_16[3];
            temp0_result_16[4] <= temp0_result_16[4];
            temp0_result_16[5] <= temp0_result_16[5];
            temp0_result_16[6] <= temp0_result_16[6];
            temp0_result_16[7] <= temp0_result_16[7];
            temp0_result_16[8] <= temp0_result_16[8];
            temp0_result_16[9] <= temp0_result_16[9];
            temp0_result_16[10] <= temp0_result_16[10];
            temp0_result_16[11] <= temp0_result_16[11];
            temp0_result_16[12] <= temp0_result_16[12];
            temp0_result_16[13] <= temp0_result_16[13];
            temp0_result_16[14] <= temp0_result_16[14];
            temp0_result_16[15] <= temp0_result_16[15];
            temp1_result_16[0] <= temp1_result_16[0];
            temp1_result_16[1] <= temp1_result_16[1];
            temp1_result_16[2] <= temp1_result_16[2];
            temp1_result_16[3] <= temp1_result_16[3];
            temp1_result_16[4] <= temp1_result_16[4];
            temp1_result_16[5] <= temp1_result_16[5];
            temp1_result_16[6] <= temp1_result_16[6];
            temp1_result_16[7] <= temp1_result_16[7];
            temp1_result_16[8] <= temp1_result_16[8];
            temp1_result_16[9] <= temp1_result_16[9];
            temp1_result_16[10] <= temp1_result_16[10];
            temp1_result_16[11] <= temp1_result_16[11];
            temp1_result_16[12] <= temp1_result_16[12];
            temp1_result_16[13] <= temp1_result_16[13];
            temp1_result_16[14] <= temp1_result_16[14];
            temp1_result_16[15] <= temp1_result_16[15];
            
            temp4_result_16[0] <= temp4_result_16[0];
            temp4_result_16[1] <= temp4_result_16[1];
            temp4_result_16[2] <= temp4_result_16[2];
            temp4_result_16[3] <= temp4_result_16[3];
            temp4_result_16[4] <= temp4_result_16[4];
            temp4_result_16[5] <= temp4_result_16[5];
            temp4_result_16[6] <= temp4_result_16[6];
            temp4_result_16[7] <= temp4_result_16[7];
            temp4_result_16[8] <= temp4_result_16[8];
            temp4_result_16[9] <= temp4_result_16[9];
            temp4_result_16[10] <= temp4_result_16[10];
            temp4_result_16[11] <= temp4_result_16[11];
            temp4_result_16[12] <= temp4_result_16[12];
            temp4_result_16[13] <= temp4_result_16[13];
            temp4_result_16[14] <= temp4_result_16[14];
            temp4_result_16[15] <= temp4_result_16[15];
            temp5_result_16[0] <= temp5_result_16[0];
            temp5_result_16[1] <= temp5_result_16[1];
            temp5_result_16[2] <= temp5_result_16[2];
            temp5_result_16[3] <= temp5_result_16[3];
            temp5_result_16[4] <= temp5_result_16[4];
            temp5_result_16[5] <= temp5_result_16[5];
            temp5_result_16[6] <= temp5_result_16[6];
            temp5_result_16[7] <= temp5_result_16[7];
            temp5_result_16[8] <= temp5_result_16[8];
            temp5_result_16[9] <= temp5_result_16[9];
            temp5_result_16[10] <= temp5_result_16[10];
            temp5_result_16[11] <= temp5_result_16[11];
            temp5_result_16[12] <= temp5_result_16[12];
            temp5_result_16[13] <= temp5_result_16[13];
            temp5_result_16[14] <= temp5_result_16[14];
            temp5_result_16[15] <= temp5_result_16[15];
            
            temp8_result_16[0] <= temp8_result_16[0];
            temp8_result_16[1] <= temp8_result_16[1];
            temp8_result_16[2] <= temp8_result_16[2];
            temp8_result_16[3] <= temp8_result_16[3];
            temp8_result_16[4] <= temp8_result_16[4];
            temp8_result_16[5] <= temp8_result_16[5];
            temp8_result_16[6] <= temp8_result_16[6];
            temp8_result_16[7] <= temp8_result_16[7];
            temp8_result_16[8] <= temp8_result_16[8];
            temp8_result_16[9] <= temp8_result_16[9];
            temp8_result_16[10] <= temp8_result_16[10];
            temp8_result_16[11] <= temp8_result_16[11];
            temp8_result_16[12] <= temp8_result_16[12];
            temp8_result_16[13] <= temp8_result_16[13];
            temp8_result_16[14] <= temp8_result_16[14];
            temp8_result_16[15] <= temp8_result_16[15];
            temp9_result_16[0] <= temp9_result_16[0];
            temp9_result_16[1] <= temp9_result_16[1];
            temp9_result_16[2] <= temp9_result_16[2];
            temp9_result_16[3] <= temp9_result_16[3];
            temp9_result_16[4] <= temp9_result_16[4];
            temp9_result_16[5] <= temp9_result_16[5];
            temp9_result_16[6] <= temp9_result_16[6];
            temp9_result_16[7] <= temp9_result_16[7];
            temp9_result_16[8] <= temp9_result_16[8];
            temp9_result_16[9] <= temp9_result_16[9];
            temp9_result_16[10] <= temp9_result_16[10];
            temp9_result_16[11] <= temp9_result_16[11];
            temp9_result_16[12] <= temp9_result_16[12];
            temp9_result_16[13] <= temp9_result_16[13];
            temp9_result_16[14] <= temp9_result_16[14];
            temp9_result_16[15] <= temp9_result_16[15];
            
            temp12_result_16[0] <= temp12_result_16[0];
            temp12_result_16[1] <= temp12_result_16[1];
            temp12_result_16[2] <= temp12_result_16[2];
            temp12_result_16[3] <= temp12_result_16[3];
            temp12_result_16[4] <= temp12_result_16[4];
            temp12_result_16[5] <= temp12_result_16[5];
            temp12_result_16[6] <= temp12_result_16[6];
            temp12_result_16[7] <= temp12_result_16[7];
            temp12_result_16[8] <= temp12_result_16[8];
            temp12_result_16[9] <= temp12_result_16[9];
            temp12_result_16[10] <= temp12_result_16[10];
            temp12_result_16[11] <= temp12_result_16[11];
            temp12_result_16[12] <= temp12_result_16[12];
            temp12_result_16[13] <= temp12_result_16[13];
            temp12_result_16[14] <= temp12_result_16[14];
            temp12_result_16[15] <= temp12_result_16[15];
            temp13_result_16[0] <= temp13_result_16[0];
            temp13_result_16[1] <= temp13_result_16[1];
            temp13_result_16[2] <= temp13_result_16[2];
            temp13_result_16[3] <= temp13_result_16[3];
            temp13_result_16[4] <= temp13_result_16[4];
            temp13_result_16[5] <= temp13_result_16[5];
            temp13_result_16[6] <= temp13_result_16[6];
            temp13_result_16[7] <= temp13_result_16[7];
            temp13_result_16[8] <= temp13_result_16[8];
            temp13_result_16[9] <= temp13_result_16[9];
            temp13_result_16[10] <= temp13_result_16[10];
            temp13_result_16[11] <= temp13_result_16[11];
            temp13_result_16[12] <= temp13_result_16[12];
            temp13_result_16[13] <= temp13_result_16[13];
            temp13_result_16[14] <= temp13_result_16[14];
            temp13_result_16[15] <= temp13_result_16[15];
            

                
            end
            endcase
        end
end

always @ (posedge clk) begin    // the state machine to add temp_result_8
        if(!rst) begin
            temp0_result_8[0] <= temp0_result_8[0];
            temp0_result_8[1] <= temp0_result_8[1];
            temp0_result_8[2] <= temp0_result_8[2];
            temp0_result_8[3] <= temp0_result_8[3];
            temp0_result_8[4] <= temp0_result_8[4];
            temp0_result_8[5] <= temp0_result_8[5];
            temp0_result_8[6] <= temp0_result_8[6];
            temp0_result_8[7] <= temp0_result_8[7];
            temp1_result_8[0] <= temp1_result_8[0];
            temp1_result_8[1] <= temp1_result_8[1];
            temp1_result_8[2] <= temp1_result_8[2];
            temp1_result_8[3] <= temp1_result_8[3];
            temp1_result_8[4] <= temp1_result_8[4];
            temp1_result_8[5] <= temp1_result_8[5];
            temp1_result_8[6] <= temp1_result_8[6];
            temp1_result_8[7] <= temp1_result_8[7];
            
            temp4_result_8[0] <= temp4_result_8[0];
            temp4_result_8[1] <= temp4_result_8[1];
            temp4_result_8[2] <= temp4_result_8[2];
            temp4_result_8[3] <= temp4_result_8[3];
            temp4_result_8[4] <= temp4_result_8[4];
            temp4_result_8[5] <= temp4_result_8[5];
            temp4_result_8[6] <= temp4_result_8[6];
            temp4_result_8[7] <= temp4_result_8[7];
            temp5_result_8[0] <= temp5_result_8[0];
            temp5_result_8[1] <= temp5_result_8[1];
            temp5_result_8[2] <= temp5_result_8[2];
            temp5_result_8[3] <= temp5_result_8[3];
            temp5_result_8[4] <= temp5_result_8[4];
            temp5_result_8[5] <= temp5_result_8[5];
            temp5_result_8[6] <= temp5_result_8[6];
            temp5_result_8[7] <= temp5_result_8[7];
            
            temp8_result_8[0] <= temp8_result_8[0];
            temp8_result_8[1] <= temp8_result_8[1];
            temp8_result_8[2] <= temp8_result_8[2];
            temp8_result_8[3] <= temp8_result_8[3];
            temp8_result_8[4] <= temp8_result_8[4];
            temp8_result_8[5] <= temp8_result_8[5];
            temp8_result_8[6] <= temp8_result_8[6];
            temp8_result_8[7] <= temp8_result_8[7];
            temp9_result_8[0] <= temp9_result_8[0];
            temp9_result_8[1] <= temp9_result_8[1];
            temp9_result_8[2] <= temp9_result_8[2];
            temp9_result_8[3] <= temp9_result_8[3];
            temp9_result_8[4] <= temp9_result_8[4];
            temp9_result_8[5] <= temp9_result_8[5];
            temp9_result_8[6] <= temp9_result_8[6];
            temp9_result_8[7] <= temp9_result_8[7];
            
            temp12_result_8[0] <= temp12_result_8[0];
            temp12_result_8[1] <= temp12_result_8[1];
            temp12_result_8[2] <= temp12_result_8[2];
            temp12_result_8[3] <= temp12_result_8[3];
            temp12_result_8[4] <= temp12_result_8[4];
            temp12_result_8[5] <= temp12_result_8[5];
            temp12_result_8[6] <= temp12_result_8[6];
            temp12_result_8[7] <= temp12_result_8[7];
            temp13_result_8[0] <= temp13_result_8[0];
            temp13_result_8[1] <= temp13_result_8[1];
            temp13_result_8[2] <= temp13_result_8[2];
            temp13_result_8[3] <= temp13_result_8[3];
            temp13_result_8[4] <= temp13_result_8[4];
            temp13_result_8[5] <= temp13_result_8[5];
            temp13_result_8[6] <= temp13_result_8[6];
            temp13_result_8[7] <= temp13_result_8[7];
            
        end
        else if (idle) begin
            temp0_result_8[0] <= temp0_result_8[0];
            temp0_result_8[1] <= temp0_result_8[1];
            temp0_result_8[2] <= temp0_result_8[2];
            temp0_result_8[3] <= temp0_result_8[3];
            temp0_result_8[4] <= temp0_result_8[4];
            temp0_result_8[5] <= temp0_result_8[5];
            temp0_result_8[6] <= temp0_result_8[6];
            temp0_result_8[7] <= temp0_result_8[7];
            temp1_result_8[0] <= temp1_result_8[0];
            temp1_result_8[1] <= temp1_result_8[1];
            temp1_result_8[2] <= temp1_result_8[2];
            temp1_result_8[3] <= temp1_result_8[3];
            temp1_result_8[4] <= temp1_result_8[4];
            temp1_result_8[5] <= temp1_result_8[5];
            temp1_result_8[6] <= temp1_result_8[6];
            temp1_result_8[7] <= temp1_result_8[7];
            
            temp4_result_8[0] <= temp4_result_8[0];
            temp4_result_8[1] <= temp4_result_8[1];
            temp4_result_8[2] <= temp4_result_8[2];
            temp4_result_8[3] <= temp4_result_8[3];
            temp4_result_8[4] <= temp4_result_8[4];
            temp4_result_8[5] <= temp4_result_8[5];
            temp4_result_8[6] <= temp4_result_8[6];
            temp4_result_8[7] <= temp4_result_8[7];
            temp5_result_8[0] <= temp5_result_8[0];
            temp5_result_8[1] <= temp5_result_8[1];
            temp5_result_8[2] <= temp5_result_8[2];
            temp5_result_8[3] <= temp5_result_8[3];
            temp5_result_8[4] <= temp5_result_8[4];
            temp5_result_8[5] <= temp5_result_8[5];
            temp5_result_8[6] <= temp5_result_8[6];
            temp5_result_8[7] <= temp5_result_8[7];
            
            temp8_result_8[0] <= temp8_result_8[0];
            temp8_result_8[1] <= temp8_result_8[1];
            temp8_result_8[2] <= temp8_result_8[2];
            temp8_result_8[3] <= temp8_result_8[3];
            temp8_result_8[4] <= temp8_result_8[4];
            temp8_result_8[5] <= temp8_result_8[5];
            temp8_result_8[6] <= temp8_result_8[6];
            temp8_result_8[7] <= temp8_result_8[7];
            temp9_result_8[0] <= temp9_result_8[0];
            temp9_result_8[1] <= temp9_result_8[1];
            temp9_result_8[2] <= temp9_result_8[2];
            temp9_result_8[3] <= temp9_result_8[3];
            temp9_result_8[4] <= temp9_result_8[4];
            temp9_result_8[5] <= temp9_result_8[5];
            temp9_result_8[6] <= temp9_result_8[6];
            temp9_result_8[7] <= temp9_result_8[7];
            
            temp12_result_8[0] <= temp12_result_8[0];
            temp12_result_8[1] <= temp12_result_8[1];
            temp12_result_8[2] <= temp12_result_8[2];
            temp12_result_8[3] <= temp12_result_8[3];
            temp12_result_8[4] <= temp12_result_8[4];
            temp12_result_8[5] <= temp12_result_8[5];
            temp12_result_8[6] <= temp12_result_8[6];
            temp12_result_8[7] <= temp12_result_8[7];
            temp13_result_8[0] <= temp13_result_8[0];
            temp13_result_8[1] <= temp13_result_8[1];
            temp13_result_8[2] <= temp13_result_8[2];
            temp13_result_8[3] <= temp13_result_8[3];
            temp13_result_8[4] <= temp13_result_8[4];
            temp13_result_8[5] <= temp13_result_8[5];
            temp13_result_8[6] <= temp13_result_8[6];
            temp13_result_8[7] <= temp13_result_8[7];
        end
        else begin
            case(state)
            Wait_Add128to64_64to32_32to16_16to8:begin
                temp0_result_8[0] <= temp0_result_16[0] + temp0_result_16[1];
                temp0_result_8[1] <= temp0_result_16[2] + temp0_result_16[3];
                temp0_result_8[2] <= temp0_result_16[4] + temp0_result_16[5];
                temp0_result_8[3] <= temp0_result_16[6] + temp0_result_16[7];
                temp0_result_8[4] <= temp0_result_16[8] + temp0_result_16[9];
                temp0_result_8[5] <= temp0_result_16[10] + temp0_result_16[11];
                temp0_result_8[6] <= temp0_result_16[12] + temp0_result_16[13];
                temp0_result_8[7] <= temp0_result_16[14] + temp0_result_16[15];
                temp1_result_8[0] <= temp1_result_16[0] + temp1_result_16[1];
                temp1_result_8[1] <= temp1_result_16[2] + temp1_result_16[3];
                temp1_result_8[2] <= temp1_result_16[4] + temp1_result_16[5];
                temp1_result_8[3] <= temp1_result_16[6] + temp1_result_16[7];
                temp1_result_8[4] <= temp1_result_16[8] + temp1_result_16[9];
                temp1_result_8[5] <= temp1_result_16[10] + temp1_result_16[11];
                temp1_result_8[6] <= temp1_result_16[12] + temp1_result_16[13];
                temp1_result_8[7] <= temp1_result_16[14] + temp1_result_16[15];
                
                temp4_result_8[0] <= temp4_result_16[0] + temp4_result_16[1];
                temp4_result_8[1] <= temp4_result_16[2] + temp4_result_16[3];
                temp4_result_8[2] <= temp4_result_16[4] + temp4_result_16[5];
                temp4_result_8[3] <= temp4_result_16[6] + temp4_result_16[7];
                temp4_result_8[4] <= temp4_result_16[8] + temp4_result_16[9];
                temp4_result_8[5] <= temp4_result_16[10] + temp4_result_16[11];
                temp4_result_8[6] <= temp4_result_16[12] + temp4_result_16[13];
                temp4_result_8[7] <= temp4_result_16[14] + temp4_result_16[15];
                temp5_result_8[0] <= temp5_result_16[0] + temp5_result_16[1];
                temp5_result_8[1] <= temp5_result_16[2] + temp5_result_16[3];
                temp5_result_8[2] <= temp5_result_16[4] + temp5_result_16[5];
                temp5_result_8[3] <= temp5_result_16[6] + temp5_result_16[7];
                temp5_result_8[4] <= temp5_result_16[8] + temp5_result_16[9];
                temp5_result_8[5] <= temp5_result_16[10] + temp5_result_16[11];
                temp5_result_8[6] <= temp5_result_16[12] + temp5_result_16[13];
                temp5_result_8[7] <= temp5_result_16[14] + temp5_result_16[15];
                
                temp8_result_8[0] <= temp8_result_16[0] + temp8_result_16[1];
                temp8_result_8[1] <= temp8_result_16[2] + temp8_result_16[3];
                temp8_result_8[2] <= temp8_result_16[4] + temp8_result_16[5];
                temp8_result_8[3] <= temp8_result_16[6] + temp8_result_16[7];
                temp8_result_8[4] <= temp8_result_16[8] + temp8_result_16[9];
                temp8_result_8[5] <= temp8_result_16[10] + temp8_result_16[11];
                temp8_result_8[6] <= temp8_result_16[12] + temp8_result_16[13];
                temp8_result_8[7] <= temp8_result_16[14] + temp8_result_16[15];
                temp9_result_8[0] <= temp9_result_16[0] + temp9_result_16[1];
                temp9_result_8[1] <= temp9_result_16[2] + temp9_result_16[3];
                temp9_result_8[2] <= temp9_result_16[4] + temp9_result_16[5];
                temp9_result_8[3] <= temp9_result_16[6] + temp9_result_16[7];
                temp9_result_8[4] <= temp9_result_16[8] + temp9_result_16[9];
                temp9_result_8[5] <= temp9_result_16[10] + temp9_result_16[11];
                temp9_result_8[6] <= temp9_result_16[12] + temp9_result_16[13];
                temp9_result_8[7] <= temp9_result_16[14] + temp9_result_16[15];
                
                temp12_result_8[0] <= temp12_result_16[0] + temp12_result_16[1];
                temp12_result_8[1] <= temp12_result_16[2] + temp12_result_16[3];
                temp12_result_8[2] <= temp12_result_16[4] + temp12_result_16[5];
                temp12_result_8[3] <= temp12_result_16[6] + temp12_result_16[7];
                temp12_result_8[4] <= temp12_result_16[8] + temp12_result_16[9];
                temp12_result_8[5] <= temp12_result_16[10] + temp12_result_16[11];
                temp12_result_8[6] <= temp12_result_16[12] + temp12_result_16[13];
                temp12_result_8[7] <= temp12_result_16[14] + temp12_result_16[15];
                temp13_result_8[0] <= temp13_result_16[0] + temp13_result_16[1];
                temp13_result_8[1] <= temp13_result_16[2] + temp13_result_16[3];
                temp13_result_8[2] <= temp13_result_16[4] + temp13_result_16[5];
                temp13_result_8[3] <= temp13_result_16[6] + temp13_result_16[7];
                temp13_result_8[4] <= temp13_result_16[8] + temp13_result_16[9];
                temp13_result_8[5] <= temp13_result_16[10] + temp13_result_16[11];
                temp13_result_8[6] <= temp13_result_16[12] + temp13_result_16[13];
                temp13_result_8[7] <= temp13_result_16[14] + temp13_result_16[15];
                

                
            end
            
            Wait_Add128to64_64to32_32to16_16to8_8to4:begin
                temp0_result_8[0] <= temp0_result_16[0] + temp0_result_16[1];
                temp0_result_8[1] <= temp0_result_16[2] + temp0_result_16[3];
                temp0_result_8[2] <= temp0_result_16[4] + temp0_result_16[5];
                temp0_result_8[3] <= temp0_result_16[6] + temp0_result_16[7];
                temp0_result_8[4] <= temp0_result_16[8] + temp0_result_16[9];
                temp0_result_8[5] <= temp0_result_16[10] + temp0_result_16[11];
                temp0_result_8[6] <= temp0_result_16[12] + temp0_result_16[13];
                temp0_result_8[7] <= temp0_result_16[14] + temp0_result_16[15];
                temp1_result_8[0] <= temp1_result_16[0] + temp1_result_16[1];
                temp1_result_8[1] <= temp1_result_16[2] + temp1_result_16[3];
                temp1_result_8[2] <= temp1_result_16[4] + temp1_result_16[5];
                temp1_result_8[3] <= temp1_result_16[6] + temp1_result_16[7];
                temp1_result_8[4] <= temp1_result_16[8] + temp1_result_16[9];
                temp1_result_8[5] <= temp1_result_16[10] + temp1_result_16[11];
                temp1_result_8[6] <= temp1_result_16[12] + temp1_result_16[13];
                temp1_result_8[7] <= temp1_result_16[14] + temp1_result_16[15];
                
                temp4_result_8[0] <= temp4_result_16[0] + temp4_result_16[1];
                temp4_result_8[1] <= temp4_result_16[2] + temp4_result_16[3];
                temp4_result_8[2] <= temp4_result_16[4] + temp4_result_16[5];
                temp4_result_8[3] <= temp4_result_16[6] + temp4_result_16[7];
                temp4_result_8[4] <= temp4_result_16[8] + temp4_result_16[9];
                temp4_result_8[5] <= temp4_result_16[10] + temp4_result_16[11];
                temp4_result_8[6] <= temp4_result_16[12] + temp4_result_16[13];
                temp4_result_8[7] <= temp4_result_16[14] + temp4_result_16[15];
                temp5_result_8[0] <= temp5_result_16[0] + temp5_result_16[1];
                temp5_result_8[1] <= temp5_result_16[2] + temp5_result_16[3];
                temp5_result_8[2] <= temp5_result_16[4] + temp5_result_16[5];
                temp5_result_8[3] <= temp5_result_16[6] + temp5_result_16[7];
                temp5_result_8[4] <= temp5_result_16[8] + temp5_result_16[9];
                temp5_result_8[5] <= temp5_result_16[10] + temp5_result_16[11];
                temp5_result_8[6] <= temp5_result_16[12] + temp5_result_16[13];
                temp5_result_8[7] <= temp5_result_16[14] + temp5_result_16[15];
                
                temp8_result_8[0] <= temp8_result_16[0] + temp8_result_16[1];
                temp8_result_8[1] <= temp8_result_16[2] + temp8_result_16[3];
                temp8_result_8[2] <= temp8_result_16[4] + temp8_result_16[5];
                temp8_result_8[3] <= temp8_result_16[6] + temp8_result_16[7];
                temp8_result_8[4] <= temp8_result_16[8] + temp8_result_16[9];
                temp8_result_8[5] <= temp8_result_16[10] + temp8_result_16[11];
                temp8_result_8[6] <= temp8_result_16[12] + temp8_result_16[13];
                temp8_result_8[7] <= temp8_result_16[14] + temp8_result_16[15];
                temp9_result_8[0] <= temp9_result_16[0] + temp9_result_16[1];
                temp9_result_8[1] <= temp9_result_16[2] + temp9_result_16[3];
                temp9_result_8[2] <= temp9_result_16[4] + temp9_result_16[5];
                temp9_result_8[3] <= temp9_result_16[6] + temp9_result_16[7];
                temp9_result_8[4] <= temp9_result_16[8] + temp9_result_16[9];
                temp9_result_8[5] <= temp9_result_16[10] + temp9_result_16[11];
                temp9_result_8[6] <= temp9_result_16[12] + temp9_result_16[13];
                temp9_result_8[7] <= temp9_result_16[14] + temp9_result_16[15];
                
                temp12_result_8[0] <= temp12_result_16[0] + temp12_result_16[1];
                temp12_result_8[1] <= temp12_result_16[2] + temp12_result_16[3];
                temp12_result_8[2] <= temp12_result_16[4] + temp12_result_16[5];
                temp12_result_8[3] <= temp12_result_16[6] + temp12_result_16[7];
                temp12_result_8[4] <= temp12_result_16[8] + temp12_result_16[9];
                temp12_result_8[5] <= temp12_result_16[10] + temp12_result_16[11];
                temp12_result_8[6] <= temp12_result_16[12] + temp12_result_16[13];
                temp12_result_8[7] <= temp12_result_16[14] + temp12_result_16[15];
                temp13_result_8[0] <= temp13_result_16[0] + temp13_result_16[1];
                temp13_result_8[1] <= temp13_result_16[2] + temp13_result_16[3];
                temp13_result_8[2] <= temp13_result_16[4] + temp13_result_16[5];
                temp13_result_8[3] <= temp13_result_16[6] + temp13_result_16[7];
                temp13_result_8[4] <= temp13_result_16[8] + temp13_result_16[9];
                temp13_result_8[5] <= temp13_result_16[10] + temp13_result_16[11];
                temp13_result_8[6] <= temp13_result_16[12] + temp13_result_16[13];
                temp13_result_8[7] <= temp13_result_16[14] + temp13_result_16[15];
            end

            Wait_Add128to64_64to32_32to16_16to8_8to4_4to2:begin
                temp0_result_8[0] <= temp0_result_16[0] + temp0_result_16[1];
                temp0_result_8[1] <= temp0_result_16[2] + temp0_result_16[3];
                temp0_result_8[2] <= temp0_result_16[4] + temp0_result_16[5];
                temp0_result_8[3] <= temp0_result_16[6] + temp0_result_16[7];
                temp0_result_8[4] <= temp0_result_16[8] + temp0_result_16[9];
                temp0_result_8[5] <= temp0_result_16[10] + temp0_result_16[11];
                temp0_result_8[6] <= temp0_result_16[12] + temp0_result_16[13];
                temp0_result_8[7] <= temp0_result_16[14] + temp0_result_16[15];
                temp1_result_8[0] <= temp1_result_16[0] + temp1_result_16[1];
                temp1_result_8[1] <= temp1_result_16[2] + temp1_result_16[3];
                temp1_result_8[2] <= temp1_result_16[4] + temp1_result_16[5];
                temp1_result_8[3] <= temp1_result_16[6] + temp1_result_16[7];
                temp1_result_8[4] <= temp1_result_16[8] + temp1_result_16[9];
                temp1_result_8[5] <= temp1_result_16[10] + temp1_result_16[11];
                temp1_result_8[6] <= temp1_result_16[12] + temp1_result_16[13];
                temp1_result_8[7] <= temp1_result_16[14] + temp1_result_16[15];
                
                temp4_result_8[0] <= temp4_result_16[0] + temp4_result_16[1];
                temp4_result_8[1] <= temp4_result_16[2] + temp4_result_16[3];
                temp4_result_8[2] <= temp4_result_16[4] + temp4_result_16[5];
                temp4_result_8[3] <= temp4_result_16[6] + temp4_result_16[7];
                temp4_result_8[4] <= temp4_result_16[8] + temp4_result_16[9];
                temp4_result_8[5] <= temp4_result_16[10] + temp4_result_16[11];
                temp4_result_8[6] <= temp4_result_16[12] + temp4_result_16[13];
                temp4_result_8[7] <= temp4_result_16[14] + temp4_result_16[15];
                temp5_result_8[0] <= temp5_result_16[0] + temp5_result_16[1];
                temp5_result_8[1] <= temp5_result_16[2] + temp5_result_16[3];
                temp5_result_8[2] <= temp5_result_16[4] + temp5_result_16[5];
                temp5_result_8[3] <= temp5_result_16[6] + temp5_result_16[7];
                temp5_result_8[4] <= temp5_result_16[8] + temp5_result_16[9];
                temp5_result_8[5] <= temp5_result_16[10] + temp5_result_16[11];
                temp5_result_8[6] <= temp5_result_16[12] + temp5_result_16[13];
                temp5_result_8[7] <= temp5_result_16[14] + temp5_result_16[15];
                
                temp8_result_8[0] <= temp8_result_16[0] + temp8_result_16[1];
                temp8_result_8[1] <= temp8_result_16[2] + temp8_result_16[3];
                temp8_result_8[2] <= temp8_result_16[4] + temp8_result_16[5];
                temp8_result_8[3] <= temp8_result_16[6] + temp8_result_16[7];
                temp8_result_8[4] <= temp8_result_16[8] + temp8_result_16[9];
                temp8_result_8[5] <= temp8_result_16[10] + temp8_result_16[11];
                temp8_result_8[6] <= temp8_result_16[12] + temp8_result_16[13];
                temp8_result_8[7] <= temp8_result_16[14] + temp8_result_16[15];
                temp9_result_8[0] <= temp9_result_16[0] + temp9_result_16[1];
                temp9_result_8[1] <= temp9_result_16[2] + temp9_result_16[3];
                temp9_result_8[2] <= temp9_result_16[4] + temp9_result_16[5];
                temp9_result_8[3] <= temp9_result_16[6] + temp9_result_16[7];
                temp9_result_8[4] <= temp9_result_16[8] + temp9_result_16[9];
                temp9_result_8[5] <= temp9_result_16[10] + temp9_result_16[11];
                temp9_result_8[6] <= temp9_result_16[12] + temp9_result_16[13];
                temp9_result_8[7] <= temp9_result_16[14] + temp9_result_16[15];
                
                temp12_result_8[0] <= temp12_result_16[0] + temp12_result_16[1];
                temp12_result_8[1] <= temp12_result_16[2] + temp12_result_16[3];
                temp12_result_8[2] <= temp12_result_16[4] + temp12_result_16[5];
                temp12_result_8[3] <= temp12_result_16[6] + temp12_result_16[7];
                temp12_result_8[4] <= temp12_result_16[8] + temp12_result_16[9];
                temp12_result_8[5] <= temp12_result_16[10] + temp12_result_16[11];
                temp12_result_8[6] <= temp12_result_16[12] + temp12_result_16[13];
                temp12_result_8[7] <= temp12_result_16[14] + temp12_result_16[15];
                temp13_result_8[0] <= temp13_result_16[0] + temp13_result_16[1];
                temp13_result_8[1] <= temp13_result_16[2] + temp13_result_16[3];
                temp13_result_8[2] <= temp13_result_16[4] + temp13_result_16[5];
                temp13_result_8[3] <= temp13_result_16[6] + temp13_result_16[7];
                temp13_result_8[4] <= temp13_result_16[8] + temp13_result_16[9];
                temp13_result_8[5] <= temp13_result_16[10] + temp13_result_16[11];
                temp13_result_8[6] <= temp13_result_16[12] + temp13_result_16[13];
                temp13_result_8[7] <= temp13_result_16[14] + temp13_result_16[15];
            end

            Wait_Add128to64_64to32_32to16_16to8_8to4_4to2_2to1:begin
                temp0_result_8[0] <= temp0_result_16[0] + temp0_result_16[1];
                temp0_result_8[1] <= temp0_result_16[2] + temp0_result_16[3];
                temp0_result_8[2] <= temp0_result_16[4] + temp0_result_16[5];
                temp0_result_8[3] <= temp0_result_16[6] + temp0_result_16[7];
                temp0_result_8[4] <= temp0_result_16[8] + temp0_result_16[9];
                temp0_result_8[5] <= temp0_result_16[10] + temp0_result_16[11];
                temp0_result_8[6] <= temp0_result_16[12] + temp0_result_16[13];
                temp0_result_8[7] <= temp0_result_16[14] + temp0_result_16[15];
                temp1_result_8[0] <= temp1_result_16[0] + temp1_result_16[1];
                temp1_result_8[1] <= temp1_result_16[2] + temp1_result_16[3];
                temp1_result_8[2] <= temp1_result_16[4] + temp1_result_16[5];
                temp1_result_8[3] <= temp1_result_16[6] + temp1_result_16[7];
                temp1_result_8[4] <= temp1_result_16[8] + temp1_result_16[9];
                temp1_result_8[5] <= temp1_result_16[10] + temp1_result_16[11];
                temp1_result_8[6] <= temp1_result_16[12] + temp1_result_16[13];
                temp1_result_8[7] <= temp1_result_16[14] + temp1_result_16[15];
                
                temp4_result_8[0] <= temp4_result_16[0] + temp4_result_16[1];
                temp4_result_8[1] <= temp4_result_16[2] + temp4_result_16[3];
                temp4_result_8[2] <= temp4_result_16[4] + temp4_result_16[5];
                temp4_result_8[3] <= temp4_result_16[6] + temp4_result_16[7];
                temp4_result_8[4] <= temp4_result_16[8] + temp4_result_16[9];
                temp4_result_8[5] <= temp4_result_16[10] + temp4_result_16[11];
                temp4_result_8[6] <= temp4_result_16[12] + temp4_result_16[13];
                temp4_result_8[7] <= temp4_result_16[14] + temp4_result_16[15];
                temp5_result_8[0] <= temp5_result_16[0] + temp5_result_16[1];
                temp5_result_8[1] <= temp5_result_16[2] + temp5_result_16[3];
                temp5_result_8[2] <= temp5_result_16[4] + temp5_result_16[5];
                temp5_result_8[3] <= temp5_result_16[6] + temp5_result_16[7];
                temp5_result_8[4] <= temp5_result_16[8] + temp5_result_16[9];
                temp5_result_8[5] <= temp5_result_16[10] + temp5_result_16[11];
                temp5_result_8[6] <= temp5_result_16[12] + temp5_result_16[13];
                temp5_result_8[7] <= temp5_result_16[14] + temp5_result_16[15];
                
                temp8_result_8[0] <= temp8_result_16[0] + temp8_result_16[1];
                temp8_result_8[1] <= temp8_result_16[2] + temp8_result_16[3];
                temp8_result_8[2] <= temp8_result_16[4] + temp8_result_16[5];
                temp8_result_8[3] <= temp8_result_16[6] + temp8_result_16[7];
                temp8_result_8[4] <= temp8_result_16[8] + temp8_result_16[9];
                temp8_result_8[5] <= temp8_result_16[10] + temp8_result_16[11];
                temp8_result_8[6] <= temp8_result_16[12] + temp8_result_16[13];
                temp8_result_8[7] <= temp8_result_16[14] + temp8_result_16[15];
                temp9_result_8[0] <= temp9_result_16[0] + temp9_result_16[1];
                temp9_result_8[1] <= temp9_result_16[2] + temp9_result_16[3];
                temp9_result_8[2] <= temp9_result_16[4] + temp9_result_16[5];
                temp9_result_8[3] <= temp9_result_16[6] + temp9_result_16[7];
                temp9_result_8[4] <= temp9_result_16[8] + temp9_result_16[9];
                temp9_result_8[5] <= temp9_result_16[10] + temp9_result_16[11];
                temp9_result_8[6] <= temp9_result_16[12] + temp9_result_16[13];
                temp9_result_8[7] <= temp9_result_16[14] + temp9_result_16[15];
                
                temp12_result_8[0] <= temp12_result_16[0] + temp12_result_16[1];
                temp12_result_8[1] <= temp12_result_16[2] + temp12_result_16[3];
                temp12_result_8[2] <= temp12_result_16[4] + temp12_result_16[5];
                temp12_result_8[3] <= temp12_result_16[6] + temp12_result_16[7];
                temp12_result_8[4] <= temp12_result_16[8] + temp12_result_16[9];
                temp12_result_8[5] <= temp12_result_16[10] + temp12_result_16[11];
                temp12_result_8[6] <= temp12_result_16[12] + temp12_result_16[13];
                temp12_result_8[7] <= temp12_result_16[14] + temp12_result_16[15];
                temp13_result_8[0] <= temp13_result_16[0] + temp13_result_16[1];
                temp13_result_8[1] <= temp13_result_16[2] + temp13_result_16[3];
                temp13_result_8[2] <= temp13_result_16[4] + temp13_result_16[5];
                temp13_result_8[3] <= temp13_result_16[6] + temp13_result_16[7];
                temp13_result_8[4] <= temp13_result_16[8] + temp13_result_16[9];
                temp13_result_8[5] <= temp13_result_16[10] + temp13_result_16[11];
                temp13_result_8[6] <= temp13_result_16[12] + temp13_result_16[13];
                temp13_result_8[7] <= temp13_result_16[14] + temp13_result_16[15];
            end
            Add128to64_64to32_32to16_16to8_8to4_4to2_2to1:begin
                temp0_result_8[0] <= temp0_result_16[0] + temp0_result_16[1];
                temp0_result_8[1] <= temp0_result_16[2] + temp0_result_16[3];
                temp0_result_8[2] <= temp0_result_16[4] + temp0_result_16[5];
                temp0_result_8[3] <= temp0_result_16[6] + temp0_result_16[7];
                temp0_result_8[4] <= temp0_result_16[8] + temp0_result_16[9];
                temp0_result_8[5] <= temp0_result_16[10] + temp0_result_16[11];
                temp0_result_8[6] <= temp0_result_16[12] + temp0_result_16[13];
                temp0_result_8[7] <= temp0_result_16[14] + temp0_result_16[15];
                temp1_result_8[0] <= temp1_result_16[0] + temp1_result_16[1];
                temp1_result_8[1] <= temp1_result_16[2] + temp1_result_16[3];
                temp1_result_8[2] <= temp1_result_16[4] + temp1_result_16[5];
                temp1_result_8[3] <= temp1_result_16[6] + temp1_result_16[7];
                temp1_result_8[4] <= temp1_result_16[8] + temp1_result_16[9];
                temp1_result_8[5] <= temp1_result_16[10] + temp1_result_16[11];
                temp1_result_8[6] <= temp1_result_16[12] + temp1_result_16[13];
                temp1_result_8[7] <= temp1_result_16[14] + temp1_result_16[15];
                
                temp4_result_8[0] <= temp4_result_16[0] + temp4_result_16[1];
                temp4_result_8[1] <= temp4_result_16[2] + temp4_result_16[3];
                temp4_result_8[2] <= temp4_result_16[4] + temp4_result_16[5];
                temp4_result_8[3] <= temp4_result_16[6] + temp4_result_16[7];
                temp4_result_8[4] <= temp4_result_16[8] + temp4_result_16[9];
                temp4_result_8[5] <= temp4_result_16[10] + temp4_result_16[11];
                temp4_result_8[6] <= temp4_result_16[12] + temp4_result_16[13];
                temp4_result_8[7] <= temp4_result_16[14] + temp4_result_16[15];
                temp5_result_8[0] <= temp5_result_16[0] + temp5_result_16[1];
                temp5_result_8[1] <= temp5_result_16[2] + temp5_result_16[3];
                temp5_result_8[2] <= temp5_result_16[4] + temp5_result_16[5];
                temp5_result_8[3] <= temp5_result_16[6] + temp5_result_16[7];
                temp5_result_8[4] <= temp5_result_16[8] + temp5_result_16[9];
                temp5_result_8[5] <= temp5_result_16[10] + temp5_result_16[11];
                temp5_result_8[6] <= temp5_result_16[12] + temp5_result_16[13];
                temp5_result_8[7] <= temp5_result_16[14] + temp5_result_16[15];
                
                temp8_result_8[0] <= temp8_result_16[0] + temp8_result_16[1];
                temp8_result_8[1] <= temp8_result_16[2] + temp8_result_16[3];
                temp8_result_8[2] <= temp8_result_16[4] + temp8_result_16[5];
                temp8_result_8[3] <= temp8_result_16[6] + temp8_result_16[7];
                temp8_result_8[4] <= temp8_result_16[8] + temp8_result_16[9];
                temp8_result_8[5] <= temp8_result_16[10] + temp8_result_16[11];
                temp8_result_8[6] <= temp8_result_16[12] + temp8_result_16[13];
                temp8_result_8[7] <= temp8_result_16[14] + temp8_result_16[15];
                temp9_result_8[0] <= temp9_result_16[0] + temp9_result_16[1];
                temp9_result_8[1] <= temp9_result_16[2] + temp9_result_16[3];
                temp9_result_8[2] <= temp9_result_16[4] + temp9_result_16[5];
                temp9_result_8[3] <= temp9_result_16[6] + temp9_result_16[7];
                temp9_result_8[4] <= temp9_result_16[8] + temp9_result_16[9];
                temp9_result_8[5] <= temp9_result_16[10] + temp9_result_16[11];
                temp9_result_8[6] <= temp9_result_16[12] + temp9_result_16[13];
                temp9_result_8[7] <= temp9_result_16[14] + temp9_result_16[15];
                
                temp12_result_8[0] <= temp12_result_16[0] + temp12_result_16[1];
                temp12_result_8[1] <= temp12_result_16[2] + temp12_result_16[3];
                temp12_result_8[2] <= temp12_result_16[4] + temp12_result_16[5];
                temp12_result_8[3] <= temp12_result_16[6] + temp12_result_16[7];
                temp12_result_8[4] <= temp12_result_16[8] + temp12_result_16[9];
                temp12_result_8[5] <= temp12_result_16[10] + temp12_result_16[11];
                temp12_result_8[6] <= temp12_result_16[12] + temp12_result_16[13];
                temp12_result_8[7] <= temp12_result_16[14] + temp12_result_16[15];
                temp13_result_8[0] <= temp13_result_16[0] + temp13_result_16[1];
                temp13_result_8[1] <= temp13_result_16[2] + temp13_result_16[3];
                temp13_result_8[2] <= temp13_result_16[4] + temp13_result_16[5];
                temp13_result_8[3] <= temp13_result_16[6] + temp13_result_16[7];
                temp13_result_8[4] <= temp13_result_16[8] + temp13_result_16[9];
                temp13_result_8[5] <= temp13_result_16[10] + temp13_result_16[11];
                temp13_result_8[6] <= temp13_result_16[12] + temp13_result_16[13];
                temp13_result_8[7] <= temp13_result_16[14] + temp13_result_16[15];
            end
            Add64to32_32to16_16to8_8to4_4to2_2to1:begin
                temp0_result_8[0] <= temp0_result_16[0] + temp0_result_16[1];
                temp0_result_8[1] <= temp0_result_16[2] + temp0_result_16[3];
                temp0_result_8[2] <= temp0_result_16[4] + temp0_result_16[5];
                temp0_result_8[3] <= temp0_result_16[6] + temp0_result_16[7];
                temp0_result_8[4] <= temp0_result_16[8] + temp0_result_16[9];
                temp0_result_8[5] <= temp0_result_16[10] + temp0_result_16[11];
                temp0_result_8[6] <= temp0_result_16[12] + temp0_result_16[13];
                temp0_result_8[7] <= temp0_result_16[14] + temp0_result_16[15];
                temp1_result_8[0] <= temp1_result_16[0] + temp1_result_16[1];
                temp1_result_8[1] <= temp1_result_16[2] + temp1_result_16[3];
                temp1_result_8[2] <= temp1_result_16[4] + temp1_result_16[5];
                temp1_result_8[3] <= temp1_result_16[6] + temp1_result_16[7];
                temp1_result_8[4] <= temp1_result_16[8] + temp1_result_16[9];
                temp1_result_8[5] <= temp1_result_16[10] + temp1_result_16[11];
                temp1_result_8[6] <= temp1_result_16[12] + temp1_result_16[13];
                temp1_result_8[7] <= temp1_result_16[14] + temp1_result_16[15];
                
                temp4_result_8[0] <= temp4_result_16[0] + temp4_result_16[1];
                temp4_result_8[1] <= temp4_result_16[2] + temp4_result_16[3];
                temp4_result_8[2] <= temp4_result_16[4] + temp4_result_16[5];
                temp4_result_8[3] <= temp4_result_16[6] + temp4_result_16[7];
                temp4_result_8[4] <= temp4_result_16[8] + temp4_result_16[9];
                temp4_result_8[5] <= temp4_result_16[10] + temp4_result_16[11];
                temp4_result_8[6] <= temp4_result_16[12] + temp4_result_16[13];
                temp4_result_8[7] <= temp4_result_16[14] + temp4_result_16[15];
                temp5_result_8[0] <= temp5_result_16[0] + temp5_result_16[1];
                temp5_result_8[1] <= temp5_result_16[2] + temp5_result_16[3];
                temp5_result_8[2] <= temp5_result_16[4] + temp5_result_16[5];
                temp5_result_8[3] <= temp5_result_16[6] + temp5_result_16[7];
                temp5_result_8[4] <= temp5_result_16[8] + temp5_result_16[9];
                temp5_result_8[5] <= temp5_result_16[10] + temp5_result_16[11];
                temp5_result_8[6] <= temp5_result_16[12] + temp5_result_16[13];
                temp5_result_8[7] <= temp5_result_16[14] + temp5_result_16[15];
                
                temp8_result_8[0] <= temp8_result_16[0] + temp8_result_16[1];
                temp8_result_8[1] <= temp8_result_16[2] + temp8_result_16[3];
                temp8_result_8[2] <= temp8_result_16[4] + temp8_result_16[5];
                temp8_result_8[3] <= temp8_result_16[6] + temp8_result_16[7];
                temp8_result_8[4] <= temp8_result_16[8] + temp8_result_16[9];
                temp8_result_8[5] <= temp8_result_16[10] + temp8_result_16[11];
                temp8_result_8[6] <= temp8_result_16[12] + temp8_result_16[13];
                temp8_result_8[7] <= temp8_result_16[14] + temp8_result_16[15];
                temp9_result_8[0] <= temp9_result_16[0] + temp9_result_16[1];
                temp9_result_8[1] <= temp9_result_16[2] + temp9_result_16[3];
                temp9_result_8[2] <= temp9_result_16[4] + temp9_result_16[5];
                temp9_result_8[3] <= temp9_result_16[6] + temp9_result_16[7];
                temp9_result_8[4] <= temp9_result_16[8] + temp9_result_16[9];
                temp9_result_8[5] <= temp9_result_16[10] + temp9_result_16[11];
                temp9_result_8[6] <= temp9_result_16[12] + temp9_result_16[13];
                temp9_result_8[7] <= temp9_result_16[14] + temp9_result_16[15];
                
                temp12_result_8[0] <= temp12_result_16[0] + temp12_result_16[1];
                temp12_result_8[1] <= temp12_result_16[2] + temp12_result_16[3];
                temp12_result_8[2] <= temp12_result_16[4] + temp12_result_16[5];
                temp12_result_8[3] <= temp12_result_16[6] + temp12_result_16[7];
                temp12_result_8[4] <= temp12_result_16[8] + temp12_result_16[9];
                temp12_result_8[5] <= temp12_result_16[10] + temp12_result_16[11];
                temp12_result_8[6] <= temp12_result_16[12] + temp12_result_16[13];
                temp12_result_8[7] <= temp12_result_16[14] + temp12_result_16[15];
                temp13_result_8[0] <= temp13_result_16[0] + temp13_result_16[1];
                temp13_result_8[1] <= temp13_result_16[2] + temp13_result_16[3];
                temp13_result_8[2] <= temp13_result_16[4] + temp13_result_16[5];
                temp13_result_8[3] <= temp13_result_16[6] + temp13_result_16[7];
                temp13_result_8[4] <= temp13_result_16[8] + temp13_result_16[9];
                temp13_result_8[5] <= temp13_result_16[10] + temp13_result_16[11];
                temp13_result_8[6] <= temp13_result_16[12] + temp13_result_16[13];
                temp13_result_8[7] <= temp13_result_16[14] + temp13_result_16[15];
            end
            Add32to16_16to8_8to4_4to2_2to1:begin
                temp0_result_8[0] <= temp0_result_16[0] + temp0_result_16[1];
                temp0_result_8[1] <= temp0_result_16[2] + temp0_result_16[3];
                temp0_result_8[2] <= temp0_result_16[4] + temp0_result_16[5];
                temp0_result_8[3] <= temp0_result_16[6] + temp0_result_16[7];
                temp0_result_8[4] <= temp0_result_16[8] + temp0_result_16[9];
                temp0_result_8[5] <= temp0_result_16[10] + temp0_result_16[11];
                temp0_result_8[6] <= temp0_result_16[12] + temp0_result_16[13];
                temp0_result_8[7] <= temp0_result_16[14] + temp0_result_16[15];
                temp1_result_8[0] <= temp1_result_16[0] + temp1_result_16[1];
                temp1_result_8[1] <= temp1_result_16[2] + temp1_result_16[3];
                temp1_result_8[2] <= temp1_result_16[4] + temp1_result_16[5];
                temp1_result_8[3] <= temp1_result_16[6] + temp1_result_16[7];
                temp1_result_8[4] <= temp1_result_16[8] + temp1_result_16[9];
                temp1_result_8[5] <= temp1_result_16[10] + temp1_result_16[11];
                temp1_result_8[6] <= temp1_result_16[12] + temp1_result_16[13];
                temp1_result_8[7] <= temp1_result_16[14] + temp1_result_16[15];
                
                temp4_result_8[0] <= temp4_result_16[0] + temp4_result_16[1];
                temp4_result_8[1] <= temp4_result_16[2] + temp4_result_16[3];
                temp4_result_8[2] <= temp4_result_16[4] + temp4_result_16[5];
                temp4_result_8[3] <= temp4_result_16[6] + temp4_result_16[7];
                temp4_result_8[4] <= temp4_result_16[8] + temp4_result_16[9];
                temp4_result_8[5] <= temp4_result_16[10] + temp4_result_16[11];
                temp4_result_8[6] <= temp4_result_16[12] + temp4_result_16[13];
                temp4_result_8[7] <= temp4_result_16[14] + temp4_result_16[15];
                temp5_result_8[0] <= temp5_result_16[0] + temp5_result_16[1];
                temp5_result_8[1] <= temp5_result_16[2] + temp5_result_16[3];
                temp5_result_8[2] <= temp5_result_16[4] + temp5_result_16[5];
                temp5_result_8[3] <= temp5_result_16[6] + temp5_result_16[7];
                temp5_result_8[4] <= temp5_result_16[8] + temp5_result_16[9];
                temp5_result_8[5] <= temp5_result_16[10] + temp5_result_16[11];
                temp5_result_8[6] <= temp5_result_16[12] + temp5_result_16[13];
                temp5_result_8[7] <= temp5_result_16[14] + temp5_result_16[15];
                
                temp8_result_8[0] <= temp8_result_16[0] + temp8_result_16[1];
                temp8_result_8[1] <= temp8_result_16[2] + temp8_result_16[3];
                temp8_result_8[2] <= temp8_result_16[4] + temp8_result_16[5];
                temp8_result_8[3] <= temp8_result_16[6] + temp8_result_16[7];
                temp8_result_8[4] <= temp8_result_16[8] + temp8_result_16[9];
                temp8_result_8[5] <= temp8_result_16[10] + temp8_result_16[11];
                temp8_result_8[6] <= temp8_result_16[12] + temp8_result_16[13];
                temp8_result_8[7] <= temp8_result_16[14] + temp8_result_16[15];
                temp9_result_8[0] <= temp9_result_16[0] + temp9_result_16[1];
                temp9_result_8[1] <= temp9_result_16[2] + temp9_result_16[3];
                temp9_result_8[2] <= temp9_result_16[4] + temp9_result_16[5];
                temp9_result_8[3] <= temp9_result_16[6] + temp9_result_16[7];
                temp9_result_8[4] <= temp9_result_16[8] + temp9_result_16[9];
                temp9_result_8[5] <= temp9_result_16[10] + temp9_result_16[11];
                temp9_result_8[6] <= temp9_result_16[12] + temp9_result_16[13];
                temp9_result_8[7] <= temp9_result_16[14] + temp9_result_16[15];
                
                temp12_result_8[0] <= temp12_result_16[0] + temp12_result_16[1];
                temp12_result_8[1] <= temp12_result_16[2] + temp12_result_16[3];
                temp12_result_8[2] <= temp12_result_16[4] + temp12_result_16[5];
                temp12_result_8[3] <= temp12_result_16[6] + temp12_result_16[7];
                temp12_result_8[4] <= temp12_result_16[8] + temp12_result_16[9];
                temp12_result_8[5] <= temp12_result_16[10] + temp12_result_16[11];
                temp12_result_8[6] <= temp12_result_16[12] + temp12_result_16[13];
                temp12_result_8[7] <= temp12_result_16[14] + temp12_result_16[15];
                temp13_result_8[0] <= temp13_result_16[0] + temp13_result_16[1];
                temp13_result_8[1] <= temp13_result_16[2] + temp13_result_16[3];
                temp13_result_8[2] <= temp13_result_16[4] + temp13_result_16[5];
                temp13_result_8[3] <= temp13_result_16[6] + temp13_result_16[7];
                temp13_result_8[4] <= temp13_result_16[8] + temp13_result_16[9];
                temp13_result_8[5] <= temp13_result_16[10] + temp13_result_16[11];
                temp13_result_8[6] <= temp13_result_16[12] + temp13_result_16[13];
                temp13_result_8[7] <= temp13_result_16[14] + temp13_result_16[15];
            end
            Add16to8_8to4_4to2_2to1:begin
                temp0_result_8[0] <= temp0_result_16[0] + temp0_result_16[1];
                temp0_result_8[1] <= temp0_result_16[2] + temp0_result_16[3];
                temp0_result_8[2] <= temp0_result_16[4] + temp0_result_16[5];
                temp0_result_8[3] <= temp0_result_16[6] + temp0_result_16[7];
                temp0_result_8[4] <= temp0_result_16[8] + temp0_result_16[9];
                temp0_result_8[5] <= temp0_result_16[10] + temp0_result_16[11];
                temp0_result_8[6] <= temp0_result_16[12] + temp0_result_16[13];
                temp0_result_8[7] <= temp0_result_16[14] + temp0_result_16[15];
                temp1_result_8[0] <= temp1_result_16[0] + temp1_result_16[1];
                temp1_result_8[1] <= temp1_result_16[2] + temp1_result_16[3];
                temp1_result_8[2] <= temp1_result_16[4] + temp1_result_16[5];
                temp1_result_8[3] <= temp1_result_16[6] + temp1_result_16[7];
                temp1_result_8[4] <= temp1_result_16[8] + temp1_result_16[9];
                temp1_result_8[5] <= temp1_result_16[10] + temp1_result_16[11];
                temp1_result_8[6] <= temp1_result_16[12] + temp1_result_16[13];
                temp1_result_8[7] <= temp1_result_16[14] + temp1_result_16[15];
                
                temp4_result_8[0] <= temp4_result_16[0] + temp4_result_16[1];
                temp4_result_8[1] <= temp4_result_16[2] + temp4_result_16[3];
                temp4_result_8[2] <= temp4_result_16[4] + temp4_result_16[5];
                temp4_result_8[3] <= temp4_result_16[6] + temp4_result_16[7];
                temp4_result_8[4] <= temp4_result_16[8] + temp4_result_16[9];
                temp4_result_8[5] <= temp4_result_16[10] + temp4_result_16[11];
                temp4_result_8[6] <= temp4_result_16[12] + temp4_result_16[13];
                temp4_result_8[7] <= temp4_result_16[14] + temp4_result_16[15];
                temp5_result_8[0] <= temp5_result_16[0] + temp5_result_16[1];
                temp5_result_8[1] <= temp5_result_16[2] + temp5_result_16[3];
                temp5_result_8[2] <= temp5_result_16[4] + temp5_result_16[5];
                temp5_result_8[3] <= temp5_result_16[6] + temp5_result_16[7];
                temp5_result_8[4] <= temp5_result_16[8] + temp5_result_16[9];
                temp5_result_8[5] <= temp5_result_16[10] + temp5_result_16[11];
                temp5_result_8[6] <= temp5_result_16[12] + temp5_result_16[13];
                temp5_result_8[7] <= temp5_result_16[14] + temp5_result_16[15];
                
                temp8_result_8[0] <= temp8_result_16[0] + temp8_result_16[1];
                temp8_result_8[1] <= temp8_result_16[2] + temp8_result_16[3];
                temp8_result_8[2] <= temp8_result_16[4] + temp8_result_16[5];
                temp8_result_8[3] <= temp8_result_16[6] + temp8_result_16[7];
                temp8_result_8[4] <= temp8_result_16[8] + temp8_result_16[9];
                temp8_result_8[5] <= temp8_result_16[10] + temp8_result_16[11];
                temp8_result_8[6] <= temp8_result_16[12] + temp8_result_16[13];
                temp8_result_8[7] <= temp8_result_16[14] + temp8_result_16[15];
                temp9_result_8[0] <= temp9_result_16[0] + temp9_result_16[1];
                temp9_result_8[1] <= temp9_result_16[2] + temp9_result_16[3];
                temp9_result_8[2] <= temp9_result_16[4] + temp9_result_16[5];
                temp9_result_8[3] <= temp9_result_16[6] + temp9_result_16[7];
                temp9_result_8[4] <= temp9_result_16[8] + temp9_result_16[9];
                temp9_result_8[5] <= temp9_result_16[10] + temp9_result_16[11];
                temp9_result_8[6] <= temp9_result_16[12] + temp9_result_16[13];
                temp9_result_8[7] <= temp9_result_16[14] + temp9_result_16[15];
                
                temp12_result_8[0] <= temp12_result_16[0] + temp12_result_16[1];
                temp12_result_8[1] <= temp12_result_16[2] + temp12_result_16[3];
                temp12_result_8[2] <= temp12_result_16[4] + temp12_result_16[5];
                temp12_result_8[3] <= temp12_result_16[6] + temp12_result_16[7];
                temp12_result_8[4] <= temp12_result_16[8] + temp12_result_16[9];
                temp12_result_8[5] <= temp12_result_16[10] + temp12_result_16[11];
                temp12_result_8[6] <= temp12_result_16[12] + temp12_result_16[13];
                temp12_result_8[7] <= temp12_result_16[14] + temp12_result_16[15];
                temp13_result_8[0] <= temp13_result_16[0] + temp13_result_16[1];
                temp13_result_8[1] <= temp13_result_16[2] + temp13_result_16[3];
                temp13_result_8[2] <= temp13_result_16[4] + temp13_result_16[5];
                temp13_result_8[3] <= temp13_result_16[6] + temp13_result_16[7];
                temp13_result_8[4] <= temp13_result_16[8] + temp13_result_16[9];
                temp13_result_8[5] <= temp13_result_16[10] + temp13_result_16[11];
                temp13_result_8[6] <= temp13_result_16[12] + temp13_result_16[13];
                temp13_result_8[7] <= temp13_result_16[14] + temp13_result_16[15];
            end
            default:begin
                temp0_result_16[0] <= temp0_result_16[0];
                temp0_result_16[1] <= temp0_result_16[1];
                temp0_result_16[2] <= temp0_result_16[2];
                temp0_result_16[3] <= temp0_result_16[3];
                temp0_result_16[4] <= temp0_result_16[4];
                temp0_result_16[5] <= temp0_result_16[5];
                temp0_result_16[6] <= temp0_result_16[6];
                temp0_result_16[7] <= temp0_result_16[7];
                temp1_result_16[0] <= temp1_result_16[0];
                temp1_result_16[1] <= temp1_result_16[1];
                temp1_result_16[2] <= temp1_result_16[2];
                temp1_result_16[3] <= temp1_result_16[3];
                temp1_result_16[4] <= temp1_result_16[4];
                temp1_result_16[5] <= temp1_result_16[5];
                temp1_result_16[6] <= temp1_result_16[6];
                temp1_result_16[7] <= temp1_result_16[7];
                
                temp4_result_16[0] <= temp4_result_16[0];
                temp4_result_16[1] <= temp4_result_16[1];
                temp4_result_16[2] <= temp4_result_16[2];
                temp4_result_16[3] <= temp4_result_16[3];
                temp4_result_16[4] <= temp4_result_16[4];
                temp4_result_16[5] <= temp4_result_16[5];
                temp4_result_16[6] <= temp4_result_16[6];
                temp4_result_16[7] <= temp4_result_16[7];
                temp5_result_16[0] <= temp5_result_16[0];
                temp5_result_16[1] <= temp5_result_16[1];
                temp5_result_16[2] <= temp5_result_16[2];
                temp5_result_16[3] <= temp5_result_16[3];
                temp5_result_16[4] <= temp5_result_16[4];
                temp5_result_16[5] <= temp5_result_16[5];
                temp5_result_16[6] <= temp5_result_16[6];
                temp5_result_16[7] <= temp5_result_16[7];
                
                temp8_result_16[0] <= temp8_result_16[0];
                temp8_result_16[1] <= temp8_result_16[1];
                temp8_result_16[2] <= temp8_result_16[2];
                temp8_result_16[3] <= temp8_result_16[3];
                temp8_result_16[4] <= temp8_result_16[4];
                temp8_result_16[5] <= temp8_result_16[5];
                temp8_result_16[6] <= temp8_result_16[6];
                temp8_result_16[7] <= temp8_result_16[7];
                temp9_result_16[0] <= temp9_result_16[0];
                temp9_result_16[1] <= temp9_result_16[1];
                temp9_result_16[2] <= temp9_result_16[2];
                temp9_result_16[3] <= temp9_result_16[3];
                temp9_result_16[4] <= temp9_result_16[4];
                temp9_result_16[5] <= temp9_result_16[5];
                temp9_result_16[6] <= temp9_result_16[6];
                temp9_result_16[7] <= temp9_result_16[7];
                
                temp12_result_16[0] <= temp12_result_16[0];
                temp12_result_16[1] <= temp12_result_16[1];
                temp12_result_16[2] <= temp12_result_16[2];
                temp12_result_16[3] <= temp12_result_16[3];
                temp12_result_16[4] <= temp12_result_16[4];
                temp12_result_16[5] <= temp12_result_16[5];
                temp12_result_16[6] <= temp12_result_16[6];
                temp12_result_16[7] <= temp12_result_16[7];
                temp13_result_16[0] <= temp13_result_16[0];
                temp13_result_16[1] <= temp13_result_16[1];
                temp13_result_16[2] <= temp13_result_16[2];
                temp13_result_16[3] <= temp13_result_16[3];
                temp13_result_16[4] <= temp13_result_16[4];
                temp13_result_16[5] <= temp13_result_16[5];
                temp13_result_16[6] <= temp13_result_16[6];
                temp13_result_16[7] <= temp13_result_16[7];
                
            end
            endcase
        end
end

always @ (posedge clk) begin    // the state machine to add temp_result_4
        if(!rst) begin
            temp0_result_4[0] <= 'd0;
            temp0_result_4[1] <= 'd0;
            temp0_result_4[2] <= 'd0;
            temp0_result_4[3] <= 'd0;
            temp1_result_4[0] <= 'd0;
            temp1_result_4[1] <= 'd0;
            temp1_result_4[2] <= 'd0;
            temp1_result_4[3] <= 'd0;
            
            temp4_result_4[0] <= 'd0;
            temp4_result_4[1] <= 'd0;
            temp4_result_4[2] <= 'd0;
            temp4_result_4[3] <= 'd0;
            temp5_result_4[0] <= 'd0;
            temp5_result_4[1] <= 'd0;
            temp5_result_4[2] <= 'd0;
            temp5_result_4[3] <= 'd0;
            
            temp8_result_4[0] <= 'd0;
            temp8_result_4[1] <= 'd0;
            temp8_result_4[2] <= 'd0;
            temp8_result_4[3] <= 'd0;
            temp9_result_4[0] <= 'd0;
            temp9_result_4[1] <= 'd0;
            temp9_result_4[2] <= 'd0;
            temp9_result_4[3] <= 'd0;
            
            temp12_result_4[0] <= 'd0;
            temp12_result_4[1] <= 'd0;
            temp12_result_4[2] <= 'd0;
            temp12_result_4[3] <= 'd0;
            temp13_result_4[0] <= 'd0;
            temp13_result_4[1] <= 'd0;
            temp13_result_4[2] <= 'd0;
            temp13_result_4[3] <= 'd0;
            
        end
        else if (idle) begin
            temp0_result_4[0] <= 'd0;
            temp0_result_4[1] <= 'd0;
            temp0_result_4[2] <= 'd0;
            temp0_result_4[3] <= 'd0;
            temp1_result_4[0] <= 'd0;
            temp1_result_4[1] <= 'd0;
            temp1_result_4[2] <= 'd0;
            temp1_result_4[3] <= 'd0;
            
            temp4_result_4[0] <= 'd0;
            temp4_result_4[1] <= 'd0;
            temp4_result_4[2] <= 'd0;
            temp4_result_4[3] <= 'd0;
            temp5_result_4[0] <= 'd0;
            temp5_result_4[1] <= 'd0;
            temp5_result_4[2] <= 'd0;
            temp5_result_4[3] <= 'd0;
            
            temp8_result_4[0] <= 'd0;
            temp8_result_4[1] <= 'd0;
            temp8_result_4[2] <= 'd0;
            temp8_result_4[3] <= 'd0;
            temp9_result_4[0] <= 'd0;
            temp9_result_4[1] <= 'd0;
            temp9_result_4[2] <= 'd0;
            temp9_result_4[3] <= 'd0;
            
            temp12_result_4[0] <= 'd0;
            temp12_result_4[1] <= 'd0;
            temp12_result_4[2] <= 'd0;
            temp12_result_4[3] <= 'd0;
            temp13_result_4[0] <= 'd0;
            temp13_result_4[1] <= 'd0;
            temp13_result_4[2] <= 'd0;
            temp13_result_4[3] <= 'd0;
        end
        else begin
            case(state)
            Wait_Add128to64_64to32_32to16_16to8_8to4:begin
                temp0_result_4[0] <= temp0_result_8[0] + temp0_result_8[1];
                temp0_result_4[1] <= temp0_result_8[2] + temp0_result_8[3];
                temp0_result_4[2] <= temp0_result_8[4] + temp0_result_8[5];
                temp0_result_4[3] <= temp0_result_8[6] + temp0_result_8[7];
                temp1_result_4[0] <= temp1_result_8[0] + temp1_result_8[1];
                temp1_result_4[1] <= temp1_result_8[2] + temp1_result_8[3];
                temp1_result_4[2] <= temp1_result_8[4] + temp1_result_8[5];
                temp1_result_4[3] <= temp1_result_8[6] + temp1_result_8[7];
                
                temp4_result_4[0] <= temp4_result_8[0] + temp4_result_8[1];
                temp4_result_4[1] <= temp4_result_8[2] + temp4_result_8[3];
                temp4_result_4[2] <= temp4_result_8[4] + temp4_result_8[5];
                temp4_result_4[3] <= temp4_result_8[6] + temp4_result_8[7];
                temp5_result_4[0] <= temp5_result_8[0] + temp5_result_8[1];
                temp5_result_4[1] <= temp5_result_8[2] + temp5_result_8[3];
                temp5_result_4[2] <= temp5_result_8[4] + temp5_result_8[5];
                temp5_result_4[3] <= temp5_result_8[6] + temp5_result_8[7];
                
                temp8_result_4[0] <= temp8_result_8[0] + temp8_result_8[1];
                temp8_result_4[1] <= temp8_result_8[2] + temp8_result_8[3];
                temp8_result_4[2] <= temp8_result_8[4] + temp8_result_8[5];
                temp8_result_4[3] <= temp8_result_8[6] + temp8_result_8[7];
                temp9_result_4[0] <= temp9_result_8[0] + temp9_result_8[1];
                temp9_result_4[1] <= temp9_result_8[2] + temp9_result_8[3];
                temp9_result_4[2] <= temp9_result_8[4] + temp9_result_8[5];
                temp9_result_4[3] <= temp9_result_8[6] + temp9_result_8[7];
                
                temp12_result_4[0] <= temp12_result_8[0] + temp12_result_8[1];
                temp12_result_4[1] <= temp12_result_8[2] + temp12_result_8[3];
                temp12_result_4[2] <= temp12_result_8[4] + temp12_result_8[5];
                temp12_result_4[3] <= temp12_result_8[6] + temp12_result_8[7];
                temp13_result_4[0] <= temp13_result_8[0] + temp13_result_8[1];
                temp13_result_4[1] <= temp13_result_8[2] + temp13_result_8[3];
                temp13_result_4[2] <= temp13_result_8[4] + temp13_result_8[5];
                temp13_result_4[3] <= temp13_result_8[6] + temp13_result_8[7];
                
            end

            Wait_Add128to64_64to32_32to16_16to8_8to4_4to2:begin
                temp0_result_4[0] <= temp0_result_8[0] + temp0_result_8[1];
                temp0_result_4[1] <= temp0_result_8[2] + temp0_result_8[3];
                temp0_result_4[2] <= temp0_result_8[4] + temp0_result_8[5];
                temp0_result_4[3] <= temp0_result_8[6] + temp0_result_8[7];
                temp1_result_4[0] <= temp1_result_8[0] + temp1_result_8[1];
                temp1_result_4[1] <= temp1_result_8[2] + temp1_result_8[3];
                temp1_result_4[2] <= temp1_result_8[4] + temp1_result_8[5];
                temp1_result_4[3] <= temp1_result_8[6] + temp1_result_8[7];
                
                temp4_result_4[0] <= temp4_result_8[0] + temp4_result_8[1];
                temp4_result_4[1] <= temp4_result_8[2] + temp4_result_8[3];
                temp4_result_4[2] <= temp4_result_8[4] + temp4_result_8[5];
                temp4_result_4[3] <= temp4_result_8[6] + temp4_result_8[7];
                temp5_result_4[0] <= temp5_result_8[0] + temp5_result_8[1];
                temp5_result_4[1] <= temp5_result_8[2] + temp5_result_8[3];
                temp5_result_4[2] <= temp5_result_8[4] + temp5_result_8[5];
                temp5_result_4[3] <= temp5_result_8[6] + temp5_result_8[7];
                
                temp8_result_4[0] <= temp8_result_8[0] + temp8_result_8[1];
                temp8_result_4[1] <= temp8_result_8[2] + temp8_result_8[3];
                temp8_result_4[2] <= temp8_result_8[4] + temp8_result_8[5];
                temp8_result_4[3] <= temp8_result_8[6] + temp8_result_8[7];
                temp9_result_4[0] <= temp9_result_8[0] + temp9_result_8[1];
                temp9_result_4[1] <= temp9_result_8[2] + temp9_result_8[3];
                temp9_result_4[2] <= temp9_result_8[4] + temp9_result_8[5];
                temp9_result_4[3] <= temp9_result_8[6] + temp9_result_8[7];
                
                temp12_result_4[0] <= temp12_result_8[0] + temp12_result_8[1];
                temp12_result_4[1] <= temp12_result_8[2] + temp12_result_8[3];
                temp12_result_4[2] <= temp12_result_8[4] + temp12_result_8[5];
                temp12_result_4[3] <= temp12_result_8[6] + temp12_result_8[7];
                temp13_result_4[0] <= temp13_result_8[0] + temp13_result_8[1];
                temp13_result_4[1] <= temp13_result_8[2] + temp13_result_8[3];
                temp13_result_4[2] <= temp13_result_8[4] + temp13_result_8[5];
                temp13_result_4[3] <= temp13_result_8[6] + temp13_result_8[7];
                
            end

            Wait_Add128to64_64to32_32to16_16to8_8to4_4to2_2to1:begin
                temp0_result_4[0] <= temp0_result_8[0] + temp0_result_8[1];
                temp0_result_4[1] <= temp0_result_8[2] + temp0_result_8[3];
                temp0_result_4[2] <= temp0_result_8[4] + temp0_result_8[5];
                temp0_result_4[3] <= temp0_result_8[6] + temp0_result_8[7];
                temp1_result_4[0] <= temp1_result_8[0] + temp1_result_8[1];
                temp1_result_4[1] <= temp1_result_8[2] + temp1_result_8[3];
                temp1_result_4[2] <= temp1_result_8[4] + temp1_result_8[5];
                temp1_result_4[3] <= temp1_result_8[6] + temp1_result_8[7];
                
                temp4_result_4[0] <= temp4_result_8[0] + temp4_result_8[1];
                temp4_result_4[1] <= temp4_result_8[2] + temp4_result_8[3];
                temp4_result_4[2] <= temp4_result_8[4] + temp4_result_8[5];
                temp4_result_4[3] <= temp4_result_8[6] + temp4_result_8[7];
                temp5_result_4[0] <= temp5_result_8[0] + temp5_result_8[1];
                temp5_result_4[1] <= temp5_result_8[2] + temp5_result_8[3];
                temp5_result_4[2] <= temp5_result_8[4] + temp5_result_8[5];
                temp5_result_4[3] <= temp5_result_8[6] + temp5_result_8[7];
                
                temp8_result_4[0] <= temp8_result_8[0] + temp8_result_8[1];
                temp8_result_4[1] <= temp8_result_8[2] + temp8_result_8[3];
                temp8_result_4[2] <= temp8_result_8[4] + temp8_result_8[5];
                temp8_result_4[3] <= temp8_result_8[6] + temp8_result_8[7];
                temp9_result_4[0] <= temp9_result_8[0] + temp9_result_8[1];
                temp9_result_4[1] <= temp9_result_8[2] + temp9_result_8[3];
                temp9_result_4[2] <= temp9_result_8[4] + temp9_result_8[5];
                temp9_result_4[3] <= temp9_result_8[6] + temp9_result_8[7];
                
                temp12_result_4[0] <= temp12_result_8[0] + temp12_result_8[1];
                temp12_result_4[1] <= temp12_result_8[2] + temp12_result_8[3];
                temp12_result_4[2] <= temp12_result_8[4] + temp12_result_8[5];
                temp12_result_4[3] <= temp12_result_8[6] + temp12_result_8[7];
                temp13_result_4[0] <= temp13_result_8[0] + temp13_result_8[1];
                temp13_result_4[1] <= temp13_result_8[2] + temp13_result_8[3];
                temp13_result_4[2] <= temp13_result_8[4] + temp13_result_8[5];
                temp13_result_4[3] <= temp13_result_8[6] + temp13_result_8[7];
                
            end
            Add128to64_64to32_32to16_16to8_8to4_4to2_2to1:begin
                temp0_result_4[0] <= temp0_result_8[0] + temp0_result_8[1];
                temp0_result_4[1] <= temp0_result_8[2] + temp0_result_8[3];
                temp0_result_4[2] <= temp0_result_8[4] + temp0_result_8[5];
                temp0_result_4[3] <= temp0_result_8[6] + temp0_result_8[7];
                temp1_result_4[0] <= temp1_result_8[0] + temp1_result_8[1];
                temp1_result_4[1] <= temp1_result_8[2] + temp1_result_8[3];
                temp1_result_4[2] <= temp1_result_8[4] + temp1_result_8[5];
                temp1_result_4[3] <= temp1_result_8[6] + temp1_result_8[7];
                
                temp4_result_4[0] <= temp4_result_8[0] + temp4_result_8[1];
                temp4_result_4[1] <= temp4_result_8[2] + temp4_result_8[3];
                temp4_result_4[2] <= temp4_result_8[4] + temp4_result_8[5];
                temp4_result_4[3] <= temp4_result_8[6] + temp4_result_8[7];
                temp5_result_4[0] <= temp5_result_8[0] + temp5_result_8[1];
                temp5_result_4[1] <= temp5_result_8[2] + temp5_result_8[3];
                temp5_result_4[2] <= temp5_result_8[4] + temp5_result_8[5];
                temp5_result_4[3] <= temp5_result_8[6] + temp5_result_8[7];
                
                temp8_result_4[0] <= temp8_result_8[0] + temp8_result_8[1];
                temp8_result_4[1] <= temp8_result_8[2] + temp8_result_8[3];
                temp8_result_4[2] <= temp8_result_8[4] + temp8_result_8[5];
                temp8_result_4[3] <= temp8_result_8[6] + temp8_result_8[7];
                temp9_result_4[0] <= temp9_result_8[0] + temp9_result_8[1];
                temp9_result_4[1] <= temp9_result_8[2] + temp9_result_8[3];
                temp9_result_4[2] <= temp9_result_8[4] + temp9_result_8[5];
                temp9_result_4[3] <= temp9_result_8[6] + temp9_result_8[7];
                
                temp12_result_4[0] <= temp12_result_8[0] + temp12_result_8[1];
                temp12_result_4[1] <= temp12_result_8[2] + temp12_result_8[3];
                temp12_result_4[2] <= temp12_result_8[4] + temp12_result_8[5];
                temp12_result_4[3] <= temp12_result_8[6] + temp12_result_8[7];
                temp13_result_4[0] <= temp13_result_8[0] + temp13_result_8[1];
                temp13_result_4[1] <= temp13_result_8[2] + temp13_result_8[3];
                temp13_result_4[2] <= temp13_result_8[4] + temp13_result_8[5];
                temp13_result_4[3] <= temp13_result_8[6] + temp13_result_8[7];
                
            end
            Add64to32_32to16_16to8_8to4_4to2_2to1:begin
                temp0_result_4[0] <= temp0_result_8[0] + temp0_result_8[1];
                temp0_result_4[1] <= temp0_result_8[2] + temp0_result_8[3];
                temp0_result_4[2] <= temp0_result_8[4] + temp0_result_8[5];
                temp0_result_4[3] <= temp0_result_8[6] + temp0_result_8[7];
                temp1_result_4[0] <= temp1_result_8[0] + temp1_result_8[1];
                temp1_result_4[1] <= temp1_result_8[2] + temp1_result_8[3];
                temp1_result_4[2] <= temp1_result_8[4] + temp1_result_8[5];
                temp1_result_4[3] <= temp1_result_8[6] + temp1_result_8[7];
                
                temp4_result_4[0] <= temp4_result_8[0] + temp4_result_8[1];
                temp4_result_4[1] <= temp4_result_8[2] + temp4_result_8[3];
                temp4_result_4[2] <= temp4_result_8[4] + temp4_result_8[5];
                temp4_result_4[3] <= temp4_result_8[6] + temp4_result_8[7];
                temp5_result_4[0] <= temp5_result_8[0] + temp5_result_8[1];
                temp5_result_4[1] <= temp5_result_8[2] + temp5_result_8[3];
                temp5_result_4[2] <= temp5_result_8[4] + temp5_result_8[5];
                temp5_result_4[3] <= temp5_result_8[6] + temp5_result_8[7];
                
                temp8_result_4[0] <= temp8_result_8[0] + temp8_result_8[1];
                temp8_result_4[1] <= temp8_result_8[2] + temp8_result_8[3];
                temp8_result_4[2] <= temp8_result_8[4] + temp8_result_8[5];
                temp8_result_4[3] <= temp8_result_8[6] + temp8_result_8[7];
                temp9_result_4[0] <= temp9_result_8[0] + temp9_result_8[1];
                temp9_result_4[1] <= temp9_result_8[2] + temp9_result_8[3];
                temp9_result_4[2] <= temp9_result_8[4] + temp9_result_8[5];
                temp9_result_4[3] <= temp9_result_8[6] + temp9_result_8[7];
                
                temp12_result_4[0] <= temp12_result_8[0] + temp12_result_8[1];
                temp12_result_4[1] <= temp12_result_8[2] + temp12_result_8[3];
                temp12_result_4[2] <= temp12_result_8[4] + temp12_result_8[5];
                temp12_result_4[3] <= temp12_result_8[6] + temp12_result_8[7];
                temp13_result_4[0] <= temp13_result_8[0] + temp13_result_8[1];
                temp13_result_4[1] <= temp13_result_8[2] + temp13_result_8[3];
                temp13_result_4[2] <= temp13_result_8[4] + temp13_result_8[5];
                temp13_result_4[3] <= temp13_result_8[6] + temp13_result_8[7];
                
            end
            Add32to16_16to8_8to4_4to2_2to1:begin
                temp0_result_4[0] <= temp0_result_8[0] + temp0_result_8[1];
                temp0_result_4[1] <= temp0_result_8[2] + temp0_result_8[3];
                temp0_result_4[2] <= temp0_result_8[4] + temp0_result_8[5];
                temp0_result_4[3] <= temp0_result_8[6] + temp0_result_8[7];
                temp1_result_4[0] <= temp1_result_8[0] + temp1_result_8[1];
                temp1_result_4[1] <= temp1_result_8[2] + temp1_result_8[3];
                temp1_result_4[2] <= temp1_result_8[4] + temp1_result_8[5];
                temp1_result_4[3] <= temp1_result_8[6] + temp1_result_8[7];
                
                temp4_result_4[0] <= temp4_result_8[0] + temp4_result_8[1];
                temp4_result_4[1] <= temp4_result_8[2] + temp4_result_8[3];
                temp4_result_4[2] <= temp4_result_8[4] + temp4_result_8[5];
                temp4_result_4[3] <= temp4_result_8[6] + temp4_result_8[7];
                temp5_result_4[0] <= temp5_result_8[0] + temp5_result_8[1];
                temp5_result_4[1] <= temp5_result_8[2] + temp5_result_8[3];
                temp5_result_4[2] <= temp5_result_8[4] + temp5_result_8[5];
                temp5_result_4[3] <= temp5_result_8[6] + temp5_result_8[7];
                
                temp8_result_4[0] <= temp8_result_8[0] + temp8_result_8[1];
                temp8_result_4[1] <= temp8_result_8[2] + temp8_result_8[3];
                temp8_result_4[2] <= temp8_result_8[4] + temp8_result_8[5];
                temp8_result_4[3] <= temp8_result_8[6] + temp8_result_8[7];
                temp9_result_4[0] <= temp9_result_8[0] + temp9_result_8[1];
                temp9_result_4[1] <= temp9_result_8[2] + temp9_result_8[3];
                temp9_result_4[2] <= temp9_result_8[4] + temp9_result_8[5];
                temp9_result_4[3] <= temp9_result_8[6] + temp9_result_8[7];
                
                temp12_result_4[0] <= temp12_result_8[0] + temp12_result_8[1];
                temp12_result_4[1] <= temp12_result_8[2] + temp12_result_8[3];
                temp12_result_4[2] <= temp12_result_8[4] + temp12_result_8[5];
                temp12_result_4[3] <= temp12_result_8[6] + temp12_result_8[7];
                temp13_result_4[0] <= temp13_result_8[0] + temp13_result_8[1];
                temp13_result_4[1] <= temp13_result_8[2] + temp13_result_8[3];
                temp13_result_4[2] <= temp13_result_8[4] + temp13_result_8[5];
                temp13_result_4[3] <= temp13_result_8[6] + temp13_result_8[7];
                
            end
            Add16to8_8to4_4to2_2to1:begin
                temp0_result_4[0] <= temp0_result_8[0] + temp0_result_8[1];
                temp0_result_4[1] <= temp0_result_8[2] + temp0_result_8[3];
                temp0_result_4[2] <= temp0_result_8[4] + temp0_result_8[5];
                temp0_result_4[3] <= temp0_result_8[6] + temp0_result_8[7];
                temp1_result_4[0] <= temp1_result_8[0] + temp1_result_8[1];
                temp1_result_4[1] <= temp1_result_8[2] + temp1_result_8[3];
                temp1_result_4[2] <= temp1_result_8[4] + temp1_result_8[5];
                temp1_result_4[3] <= temp1_result_8[6] + temp1_result_8[7];
                
                temp4_result_4[0] <= temp4_result_8[0] + temp4_result_8[1];
                temp4_result_4[1] <= temp4_result_8[2] + temp4_result_8[3];
                temp4_result_4[2] <= temp4_result_8[4] + temp4_result_8[5];
                temp4_result_4[3] <= temp4_result_8[6] + temp4_result_8[7];
                temp5_result_4[0] <= temp5_result_8[0] + temp5_result_8[1];
                temp5_result_4[1] <= temp5_result_8[2] + temp5_result_8[3];
                temp5_result_4[2] <= temp5_result_8[4] + temp5_result_8[5];
                temp5_result_4[3] <= temp5_result_8[6] + temp5_result_8[7];
                
                temp8_result_4[0] <= temp8_result_8[0] + temp8_result_8[1];
                temp8_result_4[1] <= temp8_result_8[2] + temp8_result_8[3];
                temp8_result_4[2] <= temp8_result_8[4] + temp8_result_8[5];
                temp8_result_4[3] <= temp8_result_8[6] + temp8_result_8[7];
                temp9_result_4[0] <= temp9_result_8[0] + temp9_result_8[1];
                temp9_result_4[1] <= temp9_result_8[2] + temp9_result_8[3];
                temp9_result_4[2] <= temp9_result_8[4] + temp9_result_8[5];
                temp9_result_4[3] <= temp9_result_8[6] + temp9_result_8[7];
                
                temp12_result_4[0] <= temp12_result_8[0] + temp12_result_8[1];
                temp12_result_4[1] <= temp12_result_8[2] + temp12_result_8[3];
                temp12_result_4[2] <= temp12_result_8[4] + temp12_result_8[5];
                temp12_result_4[3] <= temp12_result_8[6] + temp12_result_8[7];
                temp13_result_4[0] <= temp13_result_8[0] + temp13_result_8[1];
                temp13_result_4[1] <= temp13_result_8[2] + temp13_result_8[3];
                temp13_result_4[2] <= temp13_result_8[4] + temp13_result_8[5];
                temp13_result_4[3] <= temp13_result_8[6] + temp13_result_8[7];
                
            end
            Add8to4_4to2_2to1:begin
                temp0_result_4[0] <= temp0_result_8[0] + temp0_result_8[1];
                temp0_result_4[1] <= temp0_result_8[2] + temp0_result_8[3];
                temp0_result_4[2] <= temp0_result_8[4] + temp0_result_8[5];
                temp0_result_4[3] <= temp0_result_8[6] + temp0_result_8[7];
                temp1_result_4[0] <= temp1_result_8[0] + temp1_result_8[1];
                temp1_result_4[1] <= temp1_result_8[2] + temp1_result_8[3];
                temp1_result_4[2] <= temp1_result_8[4] + temp1_result_8[5];
                temp1_result_4[3] <= temp1_result_8[6] + temp1_result_8[7];
                
                temp4_result_4[0] <= temp4_result_8[0] + temp4_result_8[1];
                temp4_result_4[1] <= temp4_result_8[2] + temp4_result_8[3];
                temp4_result_4[2] <= temp4_result_8[4] + temp4_result_8[5];
                temp4_result_4[3] <= temp4_result_8[6] + temp4_result_8[7];
                temp5_result_4[0] <= temp5_result_8[0] + temp5_result_8[1];
                temp5_result_4[1] <= temp5_result_8[2] + temp5_result_8[3];
                temp5_result_4[2] <= temp5_result_8[4] + temp5_result_8[5];
                temp5_result_4[3] <= temp5_result_8[6] + temp5_result_8[7];
                
                temp8_result_4[0] <= temp8_result_8[0] + temp8_result_8[1];
                temp8_result_4[1] <= temp8_result_8[2] + temp8_result_8[3];
                temp8_result_4[2] <= temp8_result_8[4] + temp8_result_8[5];
                temp8_result_4[3] <= temp8_result_8[6] + temp8_result_8[7];
                temp9_result_4[0] <= temp9_result_8[0] + temp9_result_8[1];
                temp9_result_4[1] <= temp9_result_8[2] + temp9_result_8[3];
                temp9_result_4[2] <= temp9_result_8[4] + temp9_result_8[5];
                temp9_result_4[3] <= temp9_result_8[6] + temp9_result_8[7];
                
                temp12_result_4[0] <= temp12_result_8[0] + temp12_result_8[1];
                temp12_result_4[1] <= temp12_result_8[2] + temp12_result_8[3];
                temp12_result_4[2] <= temp12_result_8[4] + temp12_result_8[5];
                temp12_result_4[3] <= temp12_result_8[6] + temp12_result_8[7];
                temp13_result_4[0] <= temp13_result_8[0] + temp13_result_8[1];
                temp13_result_4[1] <= temp13_result_8[2] + temp13_result_8[3];
                temp13_result_4[2] <= temp13_result_8[4] + temp13_result_8[5];
                temp13_result_4[3] <= temp13_result_8[6] + temp13_result_8[7];
                
            end
            default:begin
                temp0_result_4[0] <= temp0_result_4[0];
                temp0_result_4[1] <= temp0_result_4[1];
                temp0_result_4[2] <= temp0_result_4[2];
                temp0_result_4[3] <= temp0_result_4[3];
                temp1_result_4[0] <= temp1_result_4[0];
                temp1_result_4[1] <= temp1_result_4[1];
                temp1_result_4[2] <= temp1_result_4[2];
                temp1_result_4[3] <= temp1_result_4[3];
                
                temp4_result_4[0] <= temp4_result_4[0];
                temp4_result_4[1] <= temp4_result_4[1];
                temp4_result_4[2] <= temp4_result_4[2];
                temp4_result_4[3] <= temp4_result_4[3];
                temp5_result_4[0] <= temp5_result_4[0];
                temp5_result_4[1] <= temp5_result_4[1];
                temp5_result_4[2] <= temp5_result_4[2];
                temp5_result_4[3] <= temp5_result_4[3];
                
                temp8_result_4[0] <= temp8_result_4[0];
                temp8_result_4[1] <= temp8_result_4[1];
                temp8_result_4[2] <= temp8_result_4[2];
                temp8_result_4[3] <= temp8_result_4[3];
                temp9_result_4[0] <= temp9_result_4[0];
                temp9_result_4[1] <= temp9_result_4[1];
                temp9_result_4[2] <= temp9_result_4[2];
                temp9_result_4[3] <= temp9_result_4[3];
                
                temp12_result_4[0] <= temp12_result_4[0];
                temp12_result_4[1] <= temp12_result_4[1];
                temp12_result_4[2] <= temp12_result_4[2];
                temp12_result_4[3] <= temp12_result_4[3];
                temp13_result_4[0] <= temp13_result_4[0];
                temp13_result_4[1] <= temp13_result_4[1];
                temp13_result_4[2] <= temp13_result_4[2];
                temp13_result_4[3] <= temp13_result_4[3];
                
            end
            endcase
        end
end


always @ (posedge clk) begin    // the state machine to add temp_result_2 and one_elements
        if(!rst) begin
            temp0_result_2[0] <= 'd0;
            temp0_result_2[1] <= 'd0;
            one_elements <= 'd0;
            temp1_result_2[0] <= 'd0;
            temp1_result_2[1] <= 'd0;
            one_elements1 <= 'd0;
            
            temp4_result_2[0] <= 'd0;
            temp4_result_2[1] <= 'd0;
            one_elements4 <= 'd0;
            temp5_result_2[0] <= 'd0;
            temp5_result_2[1] <= 'd0;
            one_elements5 <= 'd0;
            
            temp8_result_2[0] <= 'd0;
            temp8_result_2[1] <= 'd0;
            one_elements8 <= 'd0;
            temp9_result_2[0] <= 'd0;
            temp9_result_2[1] <= 'd0;
            one_elements9 <= 'd0;
            
            temp12_result_2[0] <= 'd0;
            temp12_result_2[1] <= 'd0;
            one_elements12 <= 'd0;
            temp13_result_2[0] <= 'd0;
            temp13_result_2[1] <= 'd0;
            one_elements13 <= 'd0;
            
        end
        else if (idle) begin
            temp0_result_2[0] <= 'd0;
            temp0_result_2[1] <= 'd0;
            one_elements <= 'd0;
            temp1_result_2[0] <= 'd0;
            temp1_result_2[1] <= 'd0;
            one_elements1 <= 'd0;
            
            temp4_result_2[0] <= 'd0;
            temp4_result_2[1] <= 'd0;
            one_elements4 <= 'd0;
            temp5_result_2[0] <= 'd0;
            temp5_result_2[1] <= 'd0;
            one_elements5 <= 'd0;
            
            temp8_result_2[0] <= 'd0;
            temp8_result_2[1] <= 'd0;
            one_elements8 <= 'd0;
            temp9_result_2[0] <= 'd0;
            temp9_result_2[1] <= 'd0;
            one_elements9 <= 'd0;
            
            temp12_result_2[0] <= 'd0;
            temp12_result_2[1] <= 'd0;
            one_elements12 <= 'd0;
            temp13_result_2[0] <= 'd0;
            temp13_result_2[1] <= 'd0;
            one_elements13 <= 'd0;
        end
        else begin
            case(state)
            Wait_Add128to64_64to32_32to16_16to8_8to4_4to2:begin
                temp0_result_2[0] <= temp0_result_4[0] + temp0_result_4[1];
                temp0_result_2[1] <= temp0_result_4[2] + temp0_result_4[3];
                one_elements <= one_elements;
                temp1_result_2[0] <= temp1_result_4[0] + temp1_result_4[1];
                temp1_result_2[1] <= temp1_result_4[2] + temp1_result_4[3];
                one_elements1 <= one_elements1;
                
                temp4_result_2[0] <= temp4_result_4[0] + temp4_result_4[1];
                temp4_result_2[1] <= temp4_result_4[2] + temp4_result_4[3];
                one_elements4 <= one_elements4;
                temp5_result_2[0] <= temp5_result_4[0] + temp5_result_4[1];
                temp5_result_2[1] <= temp5_result_4[2] + temp5_result_4[3];
                one_elements5 <= one_elements5;
                
                temp8_result_2[0] <= temp8_result_4[0] + temp8_result_4[1];
                temp8_result_2[1] <= temp8_result_4[2] + temp8_result_4[3];
                one_elements8 <= one_elements8;
                temp9_result_2[0] <= temp9_result_4[0] + temp9_result_4[1];
                temp9_result_2[1] <= temp9_result_4[2] + temp9_result_4[3];
                one_elements9 <= one_elements9;
                
                temp12_result_2[0] <= temp12_result_4[0] + temp12_result_4[1];
                temp12_result_2[1] <= temp12_result_4[2] + temp12_result_4[3];
                one_elements12 <= one_elements12;
                temp13_result_2[0] <= temp13_result_4[0] + temp13_result_4[1];
                temp13_result_2[1] <= temp13_result_4[2] + temp13_result_4[3];
                one_elements13 <= one_elements13;
                
            end

            Wait_Add128to64_64to32_32to16_16to8_8to4_4to2_2to1:begin
                temp0_result_2[0] <= temp0_result_4[0] + temp0_result_4[1];
                temp0_result_2[1] <= temp0_result_4[2] + temp0_result_4[3];
                one_elements <= one_elements;
                temp1_result_2[0] <= temp1_result_4[0] + temp1_result_4[1];
                temp1_result_2[1] <= temp1_result_4[2] + temp1_result_4[3];
                one_elements1 <= one_elements1;
                
                temp4_result_2[0] <= temp4_result_4[0] + temp4_result_4[1];
                temp4_result_2[1] <= temp4_result_4[2] + temp4_result_4[3];
                one_elements4 <= one_elements4;
                temp5_result_2[0] <= temp5_result_4[0] + temp5_result_4[1];
                temp5_result_2[1] <= temp5_result_4[2] + temp5_result_4[3];
                one_elements5 <= one_elements5;
                
                temp8_result_2[0] <= temp8_result_4[0] + temp8_result_4[1];
                temp8_result_2[1] <= temp8_result_4[2] + temp8_result_4[3];
                one_elements8 <= one_elements8;
                temp9_result_2[0] <= temp9_result_4[0] + temp9_result_4[1];
                temp9_result_2[1] <= temp9_result_4[2] + temp9_result_4[3];
                one_elements9 <= one_elements9;
                
                temp12_result_2[0] <= temp12_result_4[0] + temp12_result_4[1];
                temp12_result_2[1] <= temp12_result_4[2] + temp12_result_4[3];
                one_elements12 <= one_elements12;
                temp13_result_2[0] <= temp13_result_4[0] + temp13_result_4[1];
                temp13_result_2[1] <= temp13_result_4[2] + temp13_result_4[3];
                one_elements13 <= one_elements13;
            end
            Add128to64_64to32_32to16_16to8_8to4_4to2_2to1:begin
                temp0_result_2[0] <= temp0_result_4[0] + temp0_result_4[1];
                temp0_result_2[1] <= temp0_result_4[2] + temp0_result_4[3];
                one_elements <= one_elements;
                temp1_result_2[0] <= temp1_result_4[0] + temp1_result_4[1];
                temp1_result_2[1] <= temp1_result_4[2] + temp1_result_4[3];
                one_elements1 <= one_elements1;
                
                temp4_result_2[0] <= temp4_result_4[0] + temp4_result_4[1];
                temp4_result_2[1] <= temp4_result_4[2] + temp4_result_4[3];
                one_elements4 <= one_elements4;
                temp5_result_2[0] <= temp5_result_4[0] + temp5_result_4[1];
                temp5_result_2[1] <= temp5_result_4[2] + temp5_result_4[3];
                one_elements5 <= one_elements5;
                
                temp8_result_2[0] <= temp8_result_4[0] + temp8_result_4[1];
                temp8_result_2[1] <= temp8_result_4[2] + temp8_result_4[3];
                one_elements8 <= one_elements8;
                temp9_result_2[0] <= temp9_result_4[0] + temp9_result_4[1];
                temp9_result_2[1] <= temp9_result_4[2] + temp9_result_4[3];
                one_elements9 <= one_elements9;
                
                temp12_result_2[0] <= temp12_result_4[0] + temp12_result_4[1];
                temp12_result_2[1] <= temp12_result_4[2] + temp12_result_4[3];
                one_elements12 <= one_elements12;
                temp13_result_2[0] <= temp13_result_4[0] + temp13_result_4[1];
                temp13_result_2[1] <= temp13_result_4[2] + temp13_result_4[3];
                one_elements13 <= one_elements13;
            end
            Add64to32_32to16_16to8_8to4_4to2_2to1:begin
                temp0_result_2[0] <= temp0_result_4[0] + temp0_result_4[1];
                temp0_result_2[1] <= temp0_result_4[2] + temp0_result_4[3];
                one_elements <= one_elements;
                temp1_result_2[0] <= temp1_result_4[0] + temp1_result_4[1];
                temp1_result_2[1] <= temp1_result_4[2] + temp1_result_4[3];
                one_elements1 <= one_elements1;
                
                temp4_result_2[0] <= temp4_result_4[0] + temp4_result_4[1];
                temp4_result_2[1] <= temp4_result_4[2] + temp4_result_4[3];
                one_elements4 <= one_elements4;
                temp5_result_2[0] <= temp5_result_4[0] + temp5_result_4[1];
                temp5_result_2[1] <= temp5_result_4[2] + temp5_result_4[3];
                one_elements5 <= one_elements5;
                
                temp8_result_2[0] <= temp8_result_4[0] + temp8_result_4[1];
                temp8_result_2[1] <= temp8_result_4[2] + temp8_result_4[3];
                one_elements8 <= one_elements8;
                temp9_result_2[0] <= temp9_result_4[0] + temp9_result_4[1];
                temp9_result_2[1] <= temp9_result_4[2] + temp9_result_4[3];
                one_elements9 <= one_elements9;
                
                temp12_result_2[0] <= temp12_result_4[0] + temp12_result_4[1];
                temp12_result_2[1] <= temp12_result_4[2] + temp12_result_4[3];
                one_elements12 <= one_elements12;
                temp13_result_2[0] <= temp13_result_4[0] + temp13_result_4[1];
                temp13_result_2[1] <= temp13_result_4[2] + temp13_result_4[3];
                one_elements13 <= one_elements13;
            end
            Add32to16_16to8_8to4_4to2_2to1:begin
                temp0_result_2[0] <= temp0_result_4[0] + temp0_result_4[1];
                temp0_result_2[1] <= temp0_result_4[2] + temp0_result_4[3];
                one_elements <= one_elements;
                temp1_result_2[0] <= temp1_result_4[0] + temp1_result_4[1];
                temp1_result_2[1] <= temp1_result_4[2] + temp1_result_4[3];
                one_elements1 <= one_elements1;
                
                temp4_result_2[0] <= temp4_result_4[0] + temp4_result_4[1];
                temp4_result_2[1] <= temp4_result_4[2] + temp4_result_4[3];
                one_elements4 <= one_elements4;
                temp5_result_2[0] <= temp5_result_4[0] + temp5_result_4[1];
                temp5_result_2[1] <= temp5_result_4[2] + temp5_result_4[3];
                one_elements5 <= one_elements5;
                
                temp8_result_2[0] <= temp8_result_4[0] + temp8_result_4[1];
                temp8_result_2[1] <= temp8_result_4[2] + temp8_result_4[3];
                one_elements8 <= one_elements8;
                temp9_result_2[0] <= temp9_result_4[0] + temp9_result_4[1];
                temp9_result_2[1] <= temp9_result_4[2] + temp9_result_4[3];
                one_elements9 <= one_elements9;
                
                temp12_result_2[0] <= temp12_result_4[0] + temp12_result_4[1];
                temp12_result_2[1] <= temp12_result_4[2] + temp12_result_4[3];
                one_elements12 <= one_elements12;
                temp13_result_2[0] <= temp13_result_4[0] + temp13_result_4[1];
                temp13_result_2[1] <= temp13_result_4[2] + temp13_result_4[3];
                one_elements13 <= one_elements13;
            end
            Add16to8_8to4_4to2_2to1:begin
                temp0_result_2[0] <= temp0_result_4[0] + temp0_result_4[1];
                temp0_result_2[1] <= temp0_result_4[2] + temp0_result_4[3];
                one_elements <= one_elements;
                temp1_result_2[0] <= temp1_result_4[0] + temp1_result_4[1];
                temp1_result_2[1] <= temp1_result_4[2] + temp1_result_4[3];
                one_elements1 <= one_elements1;
                
                temp4_result_2[0] <= temp4_result_4[0] + temp4_result_4[1];
                temp4_result_2[1] <= temp4_result_4[2] + temp4_result_4[3];
                one_elements4 <= one_elements4;
                temp5_result_2[0] <= temp5_result_4[0] + temp5_result_4[1];
                temp5_result_2[1] <= temp5_result_4[2] + temp5_result_4[3];
                one_elements5 <= one_elements5;
                
                temp8_result_2[0] <= temp8_result_4[0] + temp8_result_4[1];
                temp8_result_2[1] <= temp8_result_4[2] + temp8_result_4[3];
                one_elements8 <= one_elements8;
                temp9_result_2[0] <= temp9_result_4[0] + temp9_result_4[1];
                temp9_result_2[1] <= temp9_result_4[2] + temp9_result_4[3];
                one_elements9 <= one_elements9;
                
                temp12_result_2[0] <= temp12_result_4[0] + temp12_result_4[1];
                temp12_result_2[1] <= temp12_result_4[2] + temp12_result_4[3];
                one_elements12 <= one_elements12;
                temp13_result_2[0] <= temp13_result_4[0] + temp13_result_4[1];
                temp13_result_2[1] <= temp13_result_4[2] + temp13_result_4[3];
                one_elements13 <= one_elements13;
            end
            Add8to4_4to2_2to1:begin
                temp0_result_2[0] <= temp0_result_4[0] + temp0_result_4[1];
                temp0_result_2[1] <= temp0_result_4[2] + temp0_result_4[3];
                one_elements <= one_elements;
                temp1_result_2[0] <= temp1_result_4[0] + temp1_result_4[1];
                temp1_result_2[1] <= temp1_result_4[2] + temp1_result_4[3];
                one_elements1 <= one_elements1;
                
                temp4_result_2[0] <= temp4_result_4[0] + temp4_result_4[1];
                temp4_result_2[1] <= temp4_result_4[2] + temp4_result_4[3];
                one_elements4 <= one_elements4;
                temp5_result_2[0] <= temp5_result_4[0] + temp5_result_4[1];
                temp5_result_2[1] <= temp5_result_4[2] + temp5_result_4[3];
                one_elements5 <= one_elements5;
                
                temp8_result_2[0] <= temp8_result_4[0] + temp8_result_4[1];
                temp8_result_2[1] <= temp8_result_4[2] + temp8_result_4[3];
                one_elements8 <= one_elements8;
                temp9_result_2[0] <= temp9_result_4[0] + temp9_result_4[1];
                temp9_result_2[1] <= temp9_result_4[2] + temp9_result_4[3];
                one_elements9 <= one_elements9;
                
                temp12_result_2[0] <= temp12_result_4[0] + temp12_result_4[1];
                temp12_result_2[1] <= temp12_result_4[2] + temp12_result_4[3];
                one_elements12 <= one_elements12;
                temp13_result_2[0] <= temp13_result_4[0] + temp13_result_4[1];
                temp13_result_2[1] <= temp13_result_4[2] + temp13_result_4[3];
                one_elements13 <= one_elements13;
            end

            Add4to2_2to1:begin
                temp0_result_2[0] <= temp0_result_4[0] + temp0_result_4[1];
                temp0_result_2[1] <= temp0_result_4[2] + temp0_result_4[3];
                one_elements <= one_elements;
                temp1_result_2[0] <= temp1_result_4[0] + temp1_result_4[1];
                temp1_result_2[1] <= temp1_result_4[2] + temp1_result_4[3];
                one_elements1 <= one_elements1;
                
                temp4_result_2[0] <= temp4_result_4[0] + temp4_result_4[1];
                temp4_result_2[1] <= temp4_result_4[2] + temp4_result_4[3];
                one_elements4 <= one_elements4;
                temp5_result_2[0] <= temp5_result_4[0] + temp5_result_4[1];
                temp5_result_2[1] <= temp5_result_4[2] + temp5_result_4[3];
                one_elements5 <= one_elements5;
                
                temp8_result_2[0] <= temp8_result_4[0] + temp8_result_4[1];
                temp8_result_2[1] <= temp8_result_4[2] + temp8_result_4[3];
                one_elements8 <= one_elements8;
                temp9_result_2[0] <= temp9_result_4[0] + temp9_result_4[1];
                temp9_result_2[1] <= temp9_result_4[2] + temp9_result_4[3];
                one_elements9 <= one_elements9;
                
                temp12_result_2[0] <= temp12_result_4[0] + temp12_result_4[1];
                temp12_result_2[1] <= temp12_result_4[2] + temp12_result_4[3];
                one_elements12 <= one_elements12;
                temp13_result_2[0] <= temp13_result_4[0] + temp13_result_4[1];
                temp13_result_2[1] <= temp13_result_4[2] + temp13_result_4[3];
                one_elements13 <= one_elements13;
            end
            Add2to1:begin
                temp0_result_2[0] <= temp0_result_2[0];
                temp0_result_2[1] <= temp0_result_2[1];
                one_elements <= temp0_result_2[0] + temp0_result_2[1];
                temp1_result_2[0] <= temp1_result_2[0];
                temp1_result_2[1] <= temp1_result_2[1];
                one_elements1 <= temp1_result_2[0] + temp1_result_2[1];
                
                temp4_result_2[0] <= temp4_result_2[0];
                temp4_result_2[1] <= temp4_result_2[1];
                one_elements4 <= temp4_result_2[0] + temp4_result_2[1];
                temp5_result_2[0] <= temp5_result_2[0];
                temp5_result_2[1] <= temp5_result_2[1];
                one_elements5 <= temp5_result_2[0] + temp5_result_2[1];
                
                temp8_result_2[0] <= temp8_result_2[0];
                temp8_result_2[1] <= temp8_result_2[1];
                one_elements8 <= temp8_result_2[0] + temp8_result_2[1];
                temp9_result_2[0] <= temp9_result_2[0];
                temp9_result_2[1] <= temp9_result_2[1];
                one_elements9 <= temp9_result_2[0] + temp9_result_2[1];
                
                temp12_result_2[0] <= temp12_result_2[0];
                temp12_result_2[1] <= temp12_result_2[1];
                one_elements12 <= temp12_result_2[0] + temp12_result_2[1];
                temp13_result_2[0] <= temp13_result_2[0];
                temp13_result_2[1] <= temp13_result_2[1];
                one_elements13 <= temp13_result_2[0] + temp13_result_2[1];
                
            end
            default:begin
                temp0_result_2[0] <= temp0_result_2[0];
                temp0_result_2[1] <= temp0_result_2[1];
                one_elements <= 'd0;
                temp1_result_2[0] <= temp1_result_2[0];
                temp1_result_2[1] <= temp1_result_2[1];
                one_elements1 <= 'd0;
                
                temp4_result_2[0] <= temp4_result_2[0];
                temp4_result_2[1] <= temp4_result_2[1];
                one_elements4 <= 'd0;
                temp5_result_2[0] <= temp5_result_2[0];
                temp5_result_2[1] <= temp5_result_2[1];
                one_elements5 <= 'd0;
                
                temp8_result_2[0] <= temp8_result_2[0];
                temp8_result_2[1] <= temp8_result_2[1];
                one_elements8 <= 'd0;
                temp9_result_2[0] <= temp9_result_2[0];
                temp9_result_2[1] <= temp9_result_2[1];
                one_elements9 <= 'd0;
                
                temp12_result_2[0] <= temp12_result_2[0];
                temp12_result_2[1] <= temp12_result_2[1];
                one_elements12 <= 'd0;
                temp13_result_2[0] <= temp13_result_2[0];
                temp13_result_2[1] <= temp13_result_2[1];
                one_elements13 <= 'd0;
                
            end
            endcase
        end
end
endmodule
